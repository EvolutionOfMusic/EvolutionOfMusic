// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.1sp1
// ALTERA_TIMESTAMP:Fri Feb  1 06:47:53 PST 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bTmxSE2QresXC8U2YgBOnIKyopPPV0unDKlKDZe8hIa4UbAn6288tM48hhwuBp/3
WRjzA9kyDwwdVn03tDfV5AlA943x+gE5P8QHzXhTBHcGCQ+PIhBLGwSP7J2d/pXm
W5x6VVJJYZ1cGAdswn/bPnCdkHB3JIQ7y+iWIb7Qmv4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16064)
BrAExLjLYnNDyLamRNUGRYt90daele05zz8/zfGcFi1zJ4aZr7ss32u6q95koxPE
ZHSoH00XB4lldDdjm4qS2LJ1x//ozv7F0b4pUJmBR4h4AiFjt81d4iDl1bURbmWr
zEXM/pWEo3Q6uqVAfN+JpoNo8u2lvCvYEROpRyutMoPEcMds3rnRsd5OX0KYzScL
q3peINI5fuyxsbn9Ay5Pa1ozn0xBJyIR5FpBvhx35YuETxtZ1kB5BJU5HxSJ6jMG
AvpFiCeljU3bRvisNgTozOiEiQ/iMz8CHpQhPA8B4AG/vpKZ5vSTv3LMLGW8jRLF
ve5qfQbO0VdbCOq4tf+6+rMiE5dH9YMN9bWBawTm3+Nv7HpaeZg0mAbAlEVkWkSQ
8TpVLwLgPru35p8PMuDmnC8cQWNCrfEda34PzHPrQZldbfAyTJU4pFLHrIMVOUMD
UlLaO8VzDSjKKUGb7C0ix9Ya5aGcn4ykz77yyYCmhRQoeSUSCJz0f2DST4cFSUjI
+cur+z0Ying6S0StKGZpz7ZPCaXf1xhwCJtU5iIgbcCydItPFFY2e/ssnnn6JpWA
ewf1+UeKRIb3sEF7lg5Gdl4EAdfpLmxPQNkVhrwqMY47ZIqiN/lkpMHnEbc68o0A
uO5LIerCS+WRwIaJ8HXb1aSS5GdO5JmOYWzPqV4hlVUhUokw/rPzDr8pF2cA9fKA
uXXLNCy7dN+0tVolZKAwRLDCwV8fukJ7yRU2KHZsYjvo7SoH8E6k74fSS60j5eaf
NU9+r8bf1opnRoZwJrgNdjbDp1oigrAR1rFVF/jawdLBeh8qxKTR8nb+kEk0ysTQ
NVK7Wh4oPGMsyfz9/kkkHXEBfuiwLwjUEU8/2Bwzh15YRRTqQLDM8jyQeSbWbvQJ
PKcuy34A6OhBZL1J0/J2L6KZ4AZ+cZomXP5h/53i4xvSvAYpLjkp9hI7sASnK1Wo
yXqxS4z0G52noZANoSmVHLsY5VHo0Xe8JsCIt+Q8j+J60WU5VffFfG+fqOuTJ/nA
rHES3f23rplPUX1PDueenHYpYSZLvZRhZwbKF0+AcnyjwJzF2XUHSYcM4f45g9E1
d7rEAygzluh797EAlYo3yD32VOEnszrUV7PeoYT1ew8K9R4GLj+jeP+WLHnjk5dw
xS2c3nXNxS4lxUiebuyyfHxAszJ5JvXJLLcWWqx0fpVMNh64nDSUG9Kvy0UQc5GR
QiF74LdiB4SM4vruiF+QVV1qFCv7ExUlPKKkw0JpCp6xDSQRkm6E2LHFNyj6jcrv
gyd5yMNfZIOKp/DJ6SXko2ta2OZvh1RGvzebDuZt3xvqIpsBiVRe7iDivpDTLaXs
TgypFEZl6Astt4u5vWT7wRwpKsoEN7xqf8Uog8kQv6QZeq1dxvh0CVJUg5sd5/QI
RGIRgJhC9pGZyRb1nHuhwS0yC2Gm5RS0hmT5fq+OH1dAjBkG4wNcf84AX63plDGm
G9Pqut+f6OEPn4jiy9TBUOhmZy2KSItvQHp5OEPiWeyKY3ejKGaalQinzexD3LUi
2Yyhtk8qQLZ5dIYW7DiK3MFcQ+5nghvCI84TdQndoY4hSzY/Yc9CUeAtio0uka6J
rSw6Q3g6aVK8aowGgUGIZ4dBbwUQt3RSg0cwDM9eHjTtHM4pGZaZvO2O+yV2dcSC
YPq4SNXLBMVsoO8npyfDvC5rlA7n3Z9hwFHz69io+7XNq4+7XyEA6+kh4bWjFsGF
Ps5seR1K/sW+4VuOMG53lf09RFdqCmekGRJgwS6N1No0KVKwvPESHtbNT7EWrPhf
NFd/HZl8RaNNBP1fnKpxFoRQWRI9RiwlaPMSV8nzwfTOMwULuplrXtkX0hvrjmID
GMV9dlhg9Gy7la4FLW4/kq9fhcTre2Ifqx8H+8Tj94uII20vPBV5bxVz6sFFpkSC
BItZHF5ASbJlu8UHJOKbg0AJzt2ds9GKPneL7BatzaUdLT/HBgCqrwx/+R7QVm+A
sTnoiToEE8p1He1oRWYYnkMynwZOMKS4PSI4VPDqfV2o+Q/KrMd0ZiqtwMx45vcZ
GUdpI1HlzB3kq/jp7nlC58xxSGWHr2G6I7HeTDvI3VPEjKz0H2K9WL+de/NCJ5TP
nIDjY4kQT/V9GVcIXlQIAWvZzrUNp2AeB3AfgpPSwIqEAoxRNAM6gDEYlVqPcmAm
a69O89JjUvOoB5NPtbhLWRHvLgE4pwVNZ7bummqcnlfI4IfyxwrZ0HqDK91tjG9w
LM1Ry8HI1RZrhRxGLkxFAsNhmMzHEwQV24H5IPS/5hj7CSaED993w5r/ZEik5KmC
LD/8ra37uEDkhX0BuvrYZTusK+MiwA58hSE44z9OPwudLvE1UoHuR1XbBse9jPNk
WYbH6UGUIk2pu+tju5kIUUm1+AAlT+s1HVmCylLrbHi5n6xtNU6sWDQDt/wDAYKc
GSA3f+6zeCZ26nr3pcDpHzBGlw/b7zGBNGszvKmun/VettcrVhRrNY7Yh3ssBDSp
CwH+ZZb91EfhIYyO5WYdQBVE3IZSfuxmIFeh4OdzUP74uozsJlvlxvxykPONDvBq
zBOmV7/KK7AYjROpmsZniF3YsfPznouYFulEazI6p2HzZl7AQWP2of8ud1mBVfPo
TDeCtZ/30hdFLOwQGE6BDKIO2suTQ6ecIHHT+Me0XVZ4ajHVTTEFdOVaKIfc8Tuv
4ECcrsNWXvjAwV/L3UmA8d5SK1myD7Gg5fThMhzI1RlrtFxdw89qHMS6L13xhSpD
gJop0yvoK8C9Z4xgQM31YD32WLRbc2RMJgY+2MJxpQ13rmXWJSzM0fHyNMcxJATm
iWPpGWgSN4vDxWEbUmefLW64em53SWCKOZd10Ydnd9eIOKZTHtQi9HlZtj7SNG6T
3TRctq0AKgb7nvFUO3ISluNrCGUxCaYaNob2kgg/F+j6DgJjzWkKzJpP8OUthkDt
CidnN1yEAWcIK1rEcXqq6DCq0v6sYwY96r6za5LCQilx5qNwGJNMmxJVyAvoVHB7
R3vKbEvK/phtJYidASwPfOqcbULS5DjEF5yrhVe+n5OBcwH1+w1FLDZt3CiFP+ob
XYYAPS006jS0gE+XmrDOA4i0UVHKEsWxt3TMOvYkFCIc7JTzUZoTq8A3K8yM1dXe
FgtqpFdPrxDbG2aV96QtPKXtes9ZmbkrtVa8+/PfN6rP4HeKv9WHO0esouIhYIu4
0ij3m/aupr/TyMyMzj4VfvRoiQKCKGo/92n+aTniDnz1in5LK/I7zeLGzlQPW7Gn
nz7RZf6yW91WW/i+uucgFfbq794u2Sl8lTkqmevwDqXWvvwDYeaHucF2I1IXtOk3
8rb4aP2gY5StfHRHe/efP4nqzX19KSnzf766UjqtmFxSoqAtz6nASKLD0ELx6+og
rxvehxcuraA3rm8GwyshbsW4uGJCLXsfK4u//Pkl4J5/32sq+7/Sfq95raGwQAVc
XbkCJ7q53ZZZRFnsQtZmpaLzMXyOQFeu/vL2TwG2eJ124qTk7ckqUYjC9V/O2XFo
E89ZcczRTfqwIqbqJOER2BWoKXOVzMRWSkJNYGGq/iiL+p00nDXmIWmWucYNuUIl
2mdclMzZJP/vmY3/wqzd8Asj86eQAT+8pdYM0nJd/wQnLA1aRBTc70hKiXw4rODq
+fIlxzi/6GLMgtZMm8bjOnn0cWtjHKULbyPg2G2dqncwuXrIRxSjZiYRtMSvxzar
B0hXnonaHqRbCuJRbPukH2j6Mab/LnyA/LxlvlaxG/z15mNuxIn9CfvQaIdH3/Lg
AopdbyHUxfJmaIk5bkWl+GAXIQiIrgtAEUY+um85iG8DqFzlwTBi+hCeQIxjWvHa
4JExZbojWfyrvbzxQd1As25wimG3h7SgudJ+jzpOT0m1tKEwV6jxbWt4pRY7MYGW
q7Ac/KdJEbkI1s8/Qz19naG6gxmse39gxiROvTQ7Bb3XX4DWwfmXUg/W8Cds+Y2/
7Gqbx6IELbrnEci2btbVeeJuNJYTeBH5y1DVtpjgl1n2a0awbf0MXupWIVxksX+e
xu82QeGVQ487NrJNb/ExD6dLkqiOMkw0IAJcMWle8MtRqHD/mF21Iu/4cwkqgLvB
nIjvHdBc/cZxfzvobSxvB6Nsct8caokoPQv9gcPdIFMn1+Muif3/YbP2gixlnLiO
Me/TDGJjdOtYMyTkHLc90WPmZuWWsVDqOLCXbaYC4/68u1R1+uZ9p/p8aPYfowTH
mL4ntWwk79VDc0tVuJWDX/KLOyVyBjV0jY69Lp2gAHW6TgyRZRFxKVdo9eSV836h
s8z/yFNHWnbcWUcHNFNt9oSYFt7YR6ty0adaKE0iUiMq3eUBMYxpvj4xyIcpdIk8
zPQrm/H3/aogROcdcSKmH51IqcysBp/kk71uY7lxAZkJqmqEvv22MlY/krzmmw8i
NLd/eeGMp6ICjS0K9EoBvItd7s9LQFffgAL9CgmCHp6QAIY1VcX+aQeazAQ0bKHX
T9Ezt8oU5Ofol1XoGS7jX1ypOOrmmYfpYsMfGZLqlUXy2ypTaFM745433BRkWM6o
RykUjEj7wKWbYCXA1ONkk0qfa7/QyqpiEdzWjUdinq1/hcjzKeomQJNJYB4XNrja
EBZDDh5UhWvU0MvLUKEu0RZZngTDPQioKt5b7/KMy11aGDrlmkHfSOg2JNDtcdJ2
McGnlT78M1JYArRC41yLGt25VVRWclBD8wHMsCrs6Bf8Hlw589pFo77Mu3d0ReeX
GnuirAfyXLmrLHX3tQjDidqnsgSjTKIG1W35+3hd3QmIG2Oe0peBTK9rVBtVGytu
XYi2tlW2ALStWdadfhBjKP+pl/RQY09rh1tnIASH6unpf8iFQAaLHeDKYpR/hQFq
9AxBpiTrFQB396YPe12HR2V0A+ZBQ3EbrsWbTvmMha0N+JGXCbHJcsO/rQHcKlag
la/2y223UiLc2uA1ebKABXYWXbebAYf9l3TuiJB4777yE36629Y9M0rIdkXtKdV9
ImbDqZwMTY3sY0OIQVlLkt8wCSfUYnushutaaELRpfeuU4HIZjC8pjYZeRvvjbTu
u5JO7oEpus98dGE3CNtcgwfrnpyiomj/38PiqW/2cgQ5bJVXY/IMSWRHaRqWW+vL
3U1Fa6VYEczBbS5oNGZxh0COAVkRUd5wEF8c6kGTauGM2tVXswHwNWygfAmMOuQg
tFZTbiAXxJMi4yARfK3upK4VScAAaI1v9zMxT758MkgmEnk6fV0k09VvCwOcfZQE
BZtIsyhq+54ICiuXoWvGr5yfsRHEROQAmnEp6p2h+i3dRWCugWtthYD8bxUe0977
EGOQ+cMVrbVx4HN6UKyQ63voQ8rJOIfasJ2vNYOS7MsoFOdTIoBTImhBJPcyQGlz
sCpNyQGVWy1pgw+BhMmC5THPPGmSgIXwaziCk+AD+zVucEgH07z/3B88WzkADd2O
X3o1F2PzIiouIfaLvMX+7oqe86PZnXSsH6GXf6QyAflIGvFtrTZtVZuHQ6/++VQe
aicUE6dp424odKSEYTummjr2FZnOjLScnvGNNctrwTO3RyMaeulSr0MsggPIs97k
p8eo22B4n7yazK5ThOj8uMlMFzbJYsIsDVjaZqJidvDYAmtLSnGG7WmDYrjK4Sjv
3ycYSkU728Bc6kfdfQrGF+fFR7MHPvpwQGQrYhkyfQM2L14A/kM3GPQMe1IluWL0
/uo7k+v+OWgmhG56hrr+ekflzONdWFpq0Q2xHbbwxXvZ5tWQyRppg7MH1V9VKTx3
2yZy+1wChr24u9AiBrsSV6Z3emRR1kczrHFyBNCWtstNhLQTn7YqFBul2y3Q9UJn
kstxDy57A9FxR94U2cRkSW7gEMZUkEWxpdtgYAL/QC2bO2mvBLnR3PxHFVNxQ6XG
Rr2QIEt6/HRkAs3yFKTib4xpYhF8T0+yErxHd7HdZBvreHSlC5Xw6XnvjHIexyoG
cIzT0zyYvHwPUtz9oum5w6TSPtbOiax94KevS/r+OHK0tPWhOZp///TZAWhamOr1
Yuze7oO8Ccx8+s9pgg2I+kNwc29qyWmrQy9AR+UpZxFRMKGaW8DJVuOEqcNWQcfK
APWhJ9nWySThKu9vD8tMRhSYimAz9YwMy4gStkoaAS9A1pwNgpFKeoEHK/mc5OOO
Ei5NBuhTyQLVL2oYr79BU0MwXHTG4g6oQDW9iSsqAKKn1SDGG0rk9EzQHhs6VVMQ
QoTnBNMhoNbmqdnR6e6gP67uyliugKl3tdnLfMeo314rQ2mH4COSBroYHVxWc8/y
LWM5qwCTz3ivdmuLmDEUwP5ZinVI5U6nHFr8C0aNm0BfB8W0dgSJghRI2YqM6EIZ
fhmb4iJKIA6EKzrPpET88ElcWKcAcZTpbj/FylH9gOdbko798X1r9/ns4B+E/WyJ
zNZOMTTjlx/zkTp6RG2AFa5Z+3g16LmvOy2A5UmTcuW2zg0wvmZvdzJbH4OmyjhW
OVVBFxNrEJ/TI3SY2gFfkpXmT1NDzirvruL9vpPvCh9a9BIhcf01DO4aNruLAaVz
ivM6f84Y0upWxDJqX+WV2M5GnRpOORu5gaHbeckeNo+rrNE1ik0tlZ8kRKJjgnKF
42M2NhT/lNm/O/rcF/pVlVoQ0rkQXyLefiEwudMH8t2Eg36a7VUu8vdIkFrjWQqG
48mebst2NFx5wFe/YbfND/tasyY0InQjNJ+QL8o5AS4YhIjxThQWDEU1GVyiOLmw
qaG3cRslTnR+9DQvy3dpozj62FTjTHMM6o4+SPw0UGzN/vZxVnx42rM3W4R6w/n1
+tHv1lKvM15DG1xQiJvKAkIbSn/+bI951WVckiFN7SZQ/0PW+0WVW5Jj5uT87385
vQHYbB47DzVn8vf0Y/tGIBPTQd5GhBBK4W0pmgc0vZ7P3B0g5cN7jNVOKK0vwsAn
siO2EshdBJqe97GPs29tzxUGeGsnFCS40Eb8ZsQ0c+RfpyR5he35hxmJP6U8E4We
bfz5P5zScNf+cvVbspy/ObloFJmF7FXOrt7XXO+eelXdpuqIuHvn/KDKlXZYoKbr
xQe9gyljY227q9jVR0j25cEIPNwP4H34lshFOnKLCDwU1Fu/OuE+bc0GW3YJJytA
1rORAz94KzrFmC66UHLcQvVdWRo4/4ws3FTwhcIUPPd2asPrl1z81dNy8u0MBwwt
/ktnlmf3MNo1IF1MM9mtXxhVt275BHBzjMyYIMjmWoybaChgYfKKjABBkJkgREbD
NYiVucf8RowO3ByBrje0sph/Vz2QPjRSqdxn0N2ReFtjMneZ9GbrDNzwH/5S9Vr4
RQ1m0IDk5pOMffxFRKseJG0OQ+hfK74MRwreLkRd9+rUMMpw3col2jr3iIaYYzWk
wfJNyaHyr9EURwMuO7VXpcTRLIVks0pggxM7zO1HjpZxujZaGxnBKFs2muJnAcYb
1oXYn7mb9RF5ajGmSuX5BmGHmk56O1KQEvGz/bpYu/0P4JYrU+T8R7aP3pOYX6BB
ZumkIUwYhcjiVlZJQ6yCMDYgxu0D5/EyrMr253tRh2hY5+tuOt91GnQexHR/dmFS
nPon/NGK6zYhoiioVRTjaK9qXxxjQZdJg6nP49yW6LXiN/2i4wUPssJmj5ULiqTW
N03n1J4ypNyn+gBzo/L17SqYw42PvKgzMmiyF+Q/9Fylj9Uq1PcH2PypjAurXTvk
rc9Ivh3GB6b7k+6xSWu1Zu7Kuf0+xd0PmBgUzHFAtYO3ZxfQNe9EgTQSIluw5g+H
jo4Tsay03yN617NCXX9L+lJlZui7ETPAaVOHr1hU/I3ZDEb87feAjP3PW5sLJQQN
vAQOSOAh5zPpglwkA5Vl3ZqjyPc/bh0greN0aup+dA0WL0P+4U1fyFBxK7Zdz1Jg
KmMdklWGJt8/IyQNCcgIpR4nmE+rflTPUGS8x6sDIFNWauCfwpcZ12vamf99p7gT
PvR5+ZDKsAQX0A03VhpemhDIUR7OErBrOohYvnESaoAErm6eYtp3/UOVTnxyW0Dc
KzCwOpNmYw81ignyLMEZokG4dsEzmhXB800BK6o66oM8X4BD1bWKjeABLaBpvW5C
IMplaNXZ3gauD0hSwX51Ei7Yl66xN/ICNhUAAWEM9UsB1q4x0ku+3L+KTBHaCCMJ
eZiYSQ3l4mvO8WPiV8GKBNGejdgkZ8jTIBMA1Xnkg2iPvYBZ5YJe46CveXCJaaQA
S8MFUimgQJ/VcRqZrF311VDtU1kKdLlj/UDi5ISvkDxV+h9TdtrpHaoV2UXxfr56
pqcZ6gCrk40E5A8aLUo1ZVpSNCxtBvCuSRhUTop8iEI6HYjIe//neecSzwotWHVJ
+X4Qpaa3Fft0RayNBfHfa+u9xbO8SWBrvnmO44azOPFgncwXQS5N+QjTjH8p2Zz/
tGe+kO6Z1ZBFoOrzzSahu6RX7408qHAzOQmuOnQw5n0Bia2ZpBWv84sga+AiGln5
ZvsMxOOkyeOwVHoNdhPEeacbJ/taHAxzLHPUjdpkR3fUaNZwnsUo4cbg9R7b0JG4
PZODNHIaChpKvgN49RgkZCv302OKa0qDTqoLXwXHPfwde+no9YOpDPIqLM4LFnXW
ZY1ay52SLB2yyTEEmsMFFFapxBUZCa0U53py/X554gB5FfVuDNL8yQiFOxs0NJSh
23zW/tA63ZRUgbuRelHBlrTQkLzN8z0zMZITS28MafGuZqjAM2Sw2v+oYdGWOjGZ
r7A27fRhDKB8PGz4bzDe1bnzPLQal9gBD1vLX3IPjGO4vi6lcd6zxzO5FIysBn7X
iqIjqVbpnPOCLYH5qrVJNsOhH4zc0AAh2Y+Gq2d5g3z7NNiROYnE9E0Evihbw/CX
LDmo2tD1BUmejzzaRsaIk19ke7yiP2+wDRObpkvWfkqYiL07XIapRVuTWOHB+jBT
CCqtaAYrmEOR3CTIFYx/+iPsbl0EbKVCYnNY+A/IevijQp3sg5b5Yd6C57o3C7sj
/WHTJn/sqbpLPJYC5uLNs3zpUbTslQyBiAuE5NAoJ/20OHoaNdaxsyesBTltB6Uw
GV8Hz+XFSpBvphgVy5In/kiLyYni9BMLo1HmRCGfGMCzPb2PoK+TOBIIPJWNkVL6
Z6UgDCRcsFPPJyrbOWgGQwb6NN35gLVczmS4gXwBRueu0xivLIhFbnw5GulrJi3k
gg/GXux/b11cMRIjMoLH00JTNtH5pP0I6z//jVwX7Z60XN+Ee/JMrqacep131nTn
qKC1p3nWWlUEjbayktCPyRTt6c2bMWJkhYNiqyW+NoYmluboFSC2W6Y9nGp90CuS
2lhTGKVwYvzv6AJ0GTHDCWRXUnMVC+Jt7eSRZ/TK6PHHh8liQxpvuP+wuY+50olf
E/amIqn9nh75uXBvywplC/B9v/rbh4QclrwLuWFVNcShd5oe+/vukFJs1p1OOXiP
vCADnfCMCvUL4HFJ3n/p6WuzxgZjAVDqPe46J9Js4QpsxMPwyWZAGmCa4dYGnIwd
FiiHdH1WkRbh66DVLrNPeOec+ZI03vqWbOdRMLJwfuuM4odCYmxt5hDqWFfcNgmE
QZOJHbiJPjQ2DwzHnZyiMHFgXwvUx8/+IAwlUZ29ELwJrADoDemU+Aq455NTqpZ7
v+bCt3BqnbyfmaTggSuGnQpQ9xILOTM0yM8+X0nBJTggfOFussFtehgMr1DgCbMN
ZYqQUbpAxIP+PYq196TcvNYKRKQG4zypbodTFvyhYzxoE8A0F01wKqcWnhVVKU54
vC/T1jnVj6sJi2RxoVAZzyqzl4osD6LZDfKTXNMr7i6NuiVj5Y1Anru9nNybn41Q
5ji8C+I//ixJKa1yPIC4oQ+f0ICmziuQo7qirilNkcNSfNxscD3S/gwuvviOT6Rj
b/nANnCLzQmzaQiEMf8NaIvNB6W8gnA7wRqpwr4fxptNhtgpNNYcocmYG4E5WaCN
Lag6XgFDzVarctTDBt62/iYGKA8O+M/wcfDFSqGkowAzApnq6jI7zN2Up02jJn5W
8CvGwGinLTcs2/IZGLC/qshRhDExeW3wxGNewUNhuBnrnHZanpoLeORQomGyduOw
CJ6QLEfmiy1ugolfYIfan6eDnrrC/A9iVu+WOUaEQSE0PD1rhsj88deTUXp1jQjN
P48P6Ab2gVhJCUUwNuk9CZHmuvpyPwmCwC888pC6aU/T34vrIpiGcBSKwK9msKNb
0YRPSLBW/D8Qoosfq8sYgpwC2m/IHTnfjg/KMoB4sqVAq0yMdOJUm8nNSxhva+kd
MuMDLgLNLBj3JWbGTgV4MJuZ22z//YnNG6WyYL96UFTIThMHlZUkBqHLLory6cRt
m7iSkQp4djZ6Rwr6Zt0KJAXPHgApdqZH5EMDWwibm1YmK9jlsQMQIiQOEjEutexk
gk0ZVfciiBF+4m66OGTZpyq+2mFJO9MKa709fASV7GYq5Mxoi09X3kO8jPuKiYVc
Wd2CSl9r/RZdNUGkcifAGsg+PDmdwBkeoKcJ4WEZZ0vJ0WjO1wIkJaICG3fGFpbk
VfSjh+6IUunPKdC0WiZ3N7VDRE7dG3pIpyr+KsoGq7uwsac7g35bJQ+LDqyAEBnI
MhrkXn687uqHgJmNNLny4eg8j/1l1C/p08+pmSXRd75LjteYSi6pFM11hAqBu6/E
gKMWEgUUbwZAfYw/06qLA3VPevpTPurSrFZz9RP5wdBXrr8ZUxjw26o2+fcDmg9R
9hhdrXxdyfSJTV8kDhOrsvC+NxdXTHh6XW5IrV63Rh9XIE/bY+FVYjcvtLk3fwPf
s9iW/qCN/Bolk1278rFO3WMyOFWLQ5ymqlqFy/DwGjY98X+F1adCaHrvCuNgeTlr
xPT8pTtOSPd6yRds0/hBEhm+V21IstnlN5wlWqd/kGmCDeUEnf+Svig9C42yU2Q1
XhpjZ5dv4pRT6St2vGISwl+8t8zee0Rjzo4AYvDtQv90ZKCLCTy21qYob8v3dZ4l
xX7RrzLK/D/PcnZbmdmF7k98Rv+ojlWN9605JI/RT473pcFWRGR7Msb4H6PfHxnD
9Liti6XycCC70dxjAgyq77tCYI2q3lX8kmqLFXn8jczAiuY5EYAhJj7uLepop2VD
HAk6GedikJ0gwFubWxxpCNz/i2FKY0uYOp/RNs8a9Qt1ZuQkEU1DKwxB4XBaA8VQ
1EtSZSWalR+qSMG3T4tGeAkgSpU+T6mKRFshhI12PJwVj3uflLa2or63H7gbkBxz
9AuLLJgZgHHmWTHJOo0H00KwZcvdDh0dXHcOYZphKfAqku4N5XyknyH8al5O0xco
XkbViL49tynuPj80LJI9I8N1AMsdGoEicp8OmB7MGigz9aCLrBTCYhFvTG6XCk8f
EzYQ16RQPLqCNUTOgjTeVNoz3OVOar1xxY9EZWse3An6REE5vcaejzx0/jCEmYCZ
viLMmWVRfBv/XFxB0QDhWzsVb5/cyIz/FsswtZSYmu9qBLUdwtGsIeloAxHPAHvJ
plo9UBi0SjO0ehI2Me76F9o+4g91yMybAOIUn7yEOvAuWTELaNN2hjMihTC1Mzju
8VlBhyc4o/W60qxpISSbF410QUkytynez1u1VvbvmRX2HNnfYu4Znv+V0RRB5GBw
p+UrBfCpQQjXqdcMZglV9Lk3wvT2pByiKtUouECjm/duJa+4eVrfp+UkZ98Pwzr5
RPp8QFn6s2XBk9YMWbVp4l0w0R1HfDUvpcjvy3ZfdenaIYLPKnHWWAg3/73N0awY
AD0Svn0C4/IyDfGPlxWvQbGwrRbFRxZhi7DqhQViD9e6f0wlpXcDU8EaYKiwQY5j
cYpYUjeMMS5mLhHBiVC1YMasCMpQcMwR/QGMlZmu+rSDN9Ll58YnhLlAFLYNBDV5
MBvkxduK0uvoFQ2q29dhYZruxSEDsXzmDHXNUK7vmsJgvqucjhq0Qzo0aUPAgaPW
TEdEnD880CymG9X7T2rWWNdjbCboNKpa0hpm59vcnqym6VBl7sxRn0cOGlhwTETh
tMR/QYzfp8TtXLbiigPyoOPj8jiP3/Bncwotl6FNp2o0LrKSXRuBZ1NsoteRjhYD
H4GHzNJZvol2ROdw1l35YWwXal3ptSa3uVNdYj17b5wvEQW019iOFKcRn5R0iPWx
8t/6pIxkdxUj+Y8GZpfylu7znskF46kWEY3gNBWchXvMK1Mu0vV2Ibiy/tgHM0Wi
QMCgFXxnvvy9p5+QDzq+sFa1bK4Pd8bBt8BxWvo2n41eg/Mz6xVNQE/+xZ1Oo7L3
1EIugKfDW5m/kRTBLM++EzwldayqHi4kWY02dtBFcRl3l5lQkeJcWqh3ZoTwA3Xp
Jd6P0YalfLKuOGSwnfcBvoos5XbefBXtMN4Q3NcfQ1F64iGVfMF7gzY4/aWiE1W7
1GUcNSaLuCycJ/wadumHgfL5r2wnIIDoXHqxOsiFHvvIVr59o7BzYo2oncT78oaS
Iv7RL8BbI+pjDXOZ7vYWQiAfvIPNdPPn1XP9qFFT5ZvGExZvBzuGuNmAFt1fl2tk
tNo6M6q5qonUj1O0F1fyIsYJiRPN3oAQrMeg/4C0gnhT7Zud8HwmLeK26ZYebW9S
7xa5dczam9z7NtQeyl/YL1dsDuqrPgGAB3ZPe3hGny6silCVMAm5ynnOE6pKC9yG
46CGw1D7tTwBsLroXUQU0934VEf7z4R9FVhfO9SbAE+oqq96GISJsSvOWQAxsQu9
hTCBnUPcQ2aW4zHXwSHOMJmleSad8fKqVac7ebrX1VoZX5VTKdW4vh6PuXlcSPNL
zguLsWdBDaaK3sasoi7CvPIoM3r5RDUuFAwrNCal1Ff+0z+1RvgJE3L9qN4HUxSG
hPs7wpE89eQTDr+OcZ7aZdw6pXk4Ls+Yr7J+SfhPI5jv7tRJMJPASx2RpRTxzFM2
DycnbB64in0ARdwOW3Xql9qxb84PWtIA1w/huoDR1Kj0J38fjQXWMxgF3xKu2FD/
+n5k37LoBwY3XILSiYDRbo7H6TL5YGQDNXE0BHjU5AfsGQYkmjJ7zEeVRmZShSri
4hkyKvMqJddcT7mG+nekbc8MNhuyVsWS+3tfXd4/XOIjZM5+unQVgtWX78SYRijJ
NAMb4xaBSDn//zvYPrCQ/JI2AEUKu1gLuvMoP8ZtNyeDMX8q+coR/hbTxXdGyvbO
nZEsFxpNcghKJkEAZ6jq3VBHRoYYjLSqbdVDonuX3waQxEp2NGGAlwlwZJOt/ix2
rbz3zIdOtS+yyPKp5xVlEf8nh+GuZgT+m05wXfOepa1Z5/gVttxy3r6dEzNlhJo5
tmODbChLJfl4Wn6SE1aU2TVCTrGxLsS/GYZLTLF6vsgyDDPRLmeFsY7e7d+z8Cqm
+1nWyGEqpemBHfnZwJGEbRjRFB5rG8zqgsNxD01138FZBXxmD6/9FFbSmn0NBvSU
xNB1krEqKu2y9lW22IX3UmLAi9wMGuS6J+7hkGEdR9w2S36++g54UV6Re8aHHzvp
MCYTlexhr+hasreoDrYxpMZKN5yOTJ4rYjkF64yuecZ7tijLGC5YGwwY6EC+Xzg2
t26ZQT4+JKlKgJfC/ZaYwIIRtqBcLWZnPF4TsbyggAhbHpu+HnOz0QeO6l/I17R9
DT5b/o7VQrywyxlSz//qYGi36mjxZ9+5v97vOldI4fpivJGuC8vjiV99q2+Fpmof
YEuaop0DbXN4OjgLoZVxK6kN/Aqhly18SxYBVZ7zDMIbqzv6wyIz+5pRRaCwVVDx
NcVx/qekbL5vilkl7WIOYjtYRNJ63OqQlvv7tOlYASKiWa1yx8F5Xk298+0v5Enh
sZWF3PsACdkM9kAn2TOpU3QyLIJEoP/NkKyMSgRwpnsyriNwIA854bI8Odco+bZy
M2NXlIq1noV2vK4JF7OT0IcrUCCX5GeraZBpFkZXOI6Wnv4K+Hfme4lG88qvGYfe
7LASsMFu8qlgl4pSKIYvnziNDU6eGb5394PgDYOq0eYZv/8zsHBW+TrRMbywS9BS
XS2/bofWYoLpiJwI+xTCnEWi6Ycxccg6cqfDE2pA5hQyR5GX94947JM3AhRccLDn
GYNOJJ+s1UMxm/iKNnoif1MbYp7BbQP7mFhShmDB0b6SQ+LiMkK6FsD12WDaE9p/
spHgOvBYKLeH9u1dRPrhRFtpiyhZUufW/4SBmCZ/u40u73LKYgDTQLnU5ACdcK5Q
1gvGggix0D2a9BK3fYNTXY8PhJFn2gVHklTYYZAKsirScRkmayei/G7kLlLVr9wS
OkZN0SyjBWmb0tRhFHJ/KHKqHfOIXZ9I02b+XYPbOmxf2BSSnaWxOtD3zxXsNl5A
wkb8Cn9z7rPl3uavo4QexyQuPHXHOkppOl62ZOcdN+oUCwPzHG8aFCM8osRT1ZEM
+Q97fQYJDvnkHLy9+KtkdYmPMEoGJ5zqquqtu/o65hWlvWL+9aB8ryrsJ0BDYVT3
T6SgHz34yFQQI7+QgXR46HyDngOsALMHXL6XO7S2+49UHDf3qL0Sh0FF5OGyDzMt
YndRa4pcK68OHL3BxvTKXztD/RTmppVomwswl9XANLuFwTd8wq0/g46FAst2xmmG
eNHses0BpkveGCY8bX3SPHGKEmEPtXYLGmU0AXeD1IaR5jCyKLtpYM8QRbgMAET0
chjI37BrSM/CJ1Xd04mft46N921K3HqUtyXrmnxDFnSg6sOEMizKJXMFs99JPMga
VLodZ3SU2PWpvx5n+sDYo4BaunQBw9Y5fROTBio92pdAtxS3JKU+jHc1T5Sp6R10
6WwYgwMAx9fq7wEEyU4IKVV5IL74BWoYwJDl5HXc4C4JOjY3B4OVR1JcW9wUetFI
+xuxPOoTZc1KYnl2+75+V2R5JzM+HGWGKl5prgk2vfHrmZ/mSi86rcbivJxtx0UJ
xIsCV3uCSjK7QkBRwtDCPwqmaqZ2mIkQDeigJGMYzJnV3mvCA+dheiIBiNjVg/eX
69ho6A9lOku1mXyg0psCfhw5fzBRUG3QX9DZoeW6Z67vxTY5JUsvW6aLR35SKcex
J5k/xZfxlupllotgRyGxRP05gAY8vEI3FcuvGLJFhMv0LI3UIUsQwzmEuaNfDMP1
lEvJ+MIWDc4oMLXxnsttai32zIlLttz8ObeD4DbklqF6smjwIDB3Fa2dPltFNcsA
SsLQu1/kIqnehCrLxGNHGRDA/3YjmeSe/Y3vzH4p6Cw+VL3gP0191b3qpwQs8P33
Am6w6hMUH14/sFdLFYLt5sxINZLYWk6t1K9eOtDo5fapPsyE7obwKz9wV1hVKJ0K
l/OLUmKIaaiVRy9NriWfX4eIg6qOdn0JvDESTRz77TsNa8cLRCUjKMi+5oBWPCPs
H9t7VMuojJTfreZpCrgyWGfOBtsEsw0itWrhsQBL16zvz1ysIaON/DKb5EcroAWc
u4YHFEg7jxJVWui3sTxgRVmMZ7880DKHv2qUJYHJ6mYYGXrhnyZjFC4txqM2f8lz
SQ8klq2xch2O5TNg3ENmzaec78ZRD/LIkNVJaflpKb6R2/1AK+r/xfMjPcx8K1Vj
KUh5OjnMYsiFf1e4uK5RT/Ie6gid6qqGEg+6/mVV5xIVE6IIHpGtieEzIASF5QtJ
nkmGbr93nF2SPjkoH7OyguWMbTgz+Yo7nKKaGQ8EXsMDOaGMSdbsVLMnj69oaEfQ
TlC7NBfNw9IUNIEReyDsgOj3+se3QmPlBNZipwjB/JMnvsF3Ft/SjMiQmluK8v+C
sVZKE2j0NsOqt1lQ8U1GKGfgcK0TdbVoKJcYjDxHu21zYRcjLGkyC1AjdXuLD9Oa
8r1gJkDiDlSwvqKTSRJl93NcDJRmHBslkVnp+EHEVnbFCaniMw1GcJM5/PrBU3EX
zbYoqsx0QK9V/tvP7e+0j2t2norlpYrbd9zFs9LrYCc9Ef+NqKYdS1oT1DYV0gY/
0n9YU5VXRzCgInqCEBC+e6KK6wCb2aOFNUROmQTHxLk9ANL596DHZ4dxiBt2lEEv
4lHpCRLplDKYG3kcsGDAC6APP8O6Nekxc6KgDYXtRN+UvlNSA9FBZgZrQED3Fe90
dLA6+pXbdSLLgWdJn6vsWZ10xsPjDHhPeX4kGuEX0tm1Y3Emed+lwPF+tGMqczMa
NBkcRJ9hSJhX3BcYIK4OFFuNbHFdB8HM0PR/MLY5kU0PtwcSecJHqW3I67w0gZbf
xj/UscaOnHpZ397GJnpy+Q+iGO5oFV4AxFsz3dPqO37/gjdEqhKy4SgSRhD6NZJc
9nnIuay5CQMud8UCJwCrV+yMdAAWoe1cWz70OMBf7m5uyKBzhs10qdGOu//1E+h3
pn6kOT3nTVFjMS5Z/PYAgCuptPZqLqX7O0P8y4HtI18fugbfwxuWPSHcMK5Kf2ov
QWD0cAdXxaCSn6lRA6fXeJCrcm3txud6dyWbzRnePwQEBvtC92j71CEcDUDbvY9e
JHNSuacrYbGnbSUElSr9Wjvj7oUsNKENaKo/1AZP9tsRT5N8Hm6/BoJ8z6SdNIKh
nKzfv0Pqvijcth7By5IyDz0IFNfTMwZBzXstY2C2xLypwfJlHXvCy4EQcLGpi8WL
0pKAnJi6CJa7HB0xKRVBZR6Y2QcAIOq8+gh4J8gEE/9sDyTu0JlYWq6ZuTRvr7kt
BBvpOVRVIBatNaZ5puZLHLE+jCP/TtPr8wv82VonlU0PhaIhsCSYlqUifBLTxtj3
GuYIBm9ymxSofiuS1nH4Uuy6l4RaQfissFoGLGsDYN8MW5G5xdAbSVYDdWWDxHwD
/4Wz0bub1ih6dP4HutOIR8fhrYY83w49n+ao6aF6o0dc9JdJYnUaYDVlWRJv/XNx
C/J9J4a3vgmRf/EHlr04+HTPgELcQYCD/iCMju1/BScsnNTFiwibB5VxSURzyCiD
nT9gLMmZEKHY2xfFTwPJqegdtKmq+rkGlRPxg/V/uIIBfMPiVuphMQwPB7Ft2RoR
4Lqqm3qL7EiRbe+EA9m8NwLTI1ToA+YerTAQSvMZPDJU7ZLDnujBETwHKrYVShTx
A5aSnsO9MbfU+EwrwrvIg4wuh8plEC2ZhpNetww5IzXzK1pEUflDIwS6ADh0weZQ
r6Ec9VRrasI+rH6MZABJNB5auxyFFupUdc65Lxqe5iaLodLO+AWFEhlS0Ngl0zvj
Dg0GeQzoz85D02DdRg+hdRO0xl0T7lff2+xyjws45uZRr3VruwCWn6I1GjVcE/17
tep22taxqi7d63n7YYRAbqF7E38Ui++c4mLhaGb5N72/0lBOdhYuaDGOWGqXLX0g
FUu0HgNjuYkFmD/8ehfmlDyD2L/fl60xPTdQOZLI3rOygIsnCdZfomNpOFvEU1+s
8O9utLJLXnCWFoYpjiHfYte16ykfNAqgKxDTFSo3jYBQegQzyn6hzdTxeG8pMSQP
ppyskLO+F4DG2+FBMCctVHIJ4sIjdr85fxUFVpJbzaJg8lehgillF2km5TS/jM7k
G2W+UDE3cZHfKeEP2vizVc+wLQvKmVaHrjvdyL5xeGC82WrP2Ja4oUQDzKDMkwXu
WAZuUCRRp/Us6Q46C8RKC1KLthCDZBi8d6bXhDh1+dza1fhY0LD9NigNWsiREJLt
BP/bLSUJYn2yKs943MgbEviRDXQ9wYXvHrwU2q7tJ4EKyTKH3ij6xEQ/hZNTtZ7e
+D5VA/OgMC0FjVDmgIhKWu7NO4DN7Yx5aEl3JVJxUHR8fcnPN9zAIt5rYqm48wVc
BvvlwCdXT5I4Y9xe5at77XHgdFn092TPzm1mqoMIpVkQqvW7l+vhJI8+V2xUGic1
Npf5HHZ2mUPkysdIAftDI2rGQuP+Q/Ao6zKdv4mwgkI/9H2Igt0pDqu4UH/Ht0pv
Pt+gM4qWuwsoNWuRT4u/BgAuEa46zQttL+8CtEDYzbN72ehXkPfQFX+CuW8tw23/
jnnn4/KHzjxSgV/5Hon6iCEqO/eZ/h+EV3LN3i+SYQdCRtx6L9ICuxz0uBSPMIxW
J9crNcOoGxpqyuU5WSZ5jbSDFgUs2TFLOMfilmEHsUb5thGVQqQZfcKwa9cOPMC0
u+5IVxBnG8t09XA4opGXvHFDNb0sS+XT7pFp84idPB5R7khHUopBBE6ypAnUFuW0
+k9uvsmYUkNrLp9umcd9x2GzmEAsB/hy3DAGdrxCSpNSpD36axF3UKXnnoKmyx11
BJJeoVHF7SzSwtBDQQMcmVOQcnkglF4bo4BpmiG0v1Cama2rvzDaHoFXn+zCVm7L
UDtmdqgNBGWs06aMQIG8ybtw/Od7E7N3S8itjf2ROs3oE2xHVpciEG/mwEXSvku1
Q2SIQyFmGZGspPOd60Cp/TLBpFeW43q2gbJ0FmYun9yzWxJ0ukYLqymHIOFEzPkx
BwHL/SzYAiC19h+oi8OAfq49H47qjr7xi4vSgTk1JopyuLOXrG2ye3BI1tRhCkbJ
c2lnyaFfiVg8m714RCyKfRIQ1sUn9l03zX0MbfF1LEMcTEwq6hS8kTE1qIcW3/g4
MbnYzHpa/+FJyjC4oLwuGVfXCl1bKcNVDg00rNEeKDOGBYPE+54v6BRmMAtzAzJF
BG2qzxQiRLJIKbnfC6smuA8nGvutrkuG2GoC+1pZY7WzUBGAWHl2QtxPdJjUKTx1
Q847Q+pKMMRVRfXK+/bkD8836N3I+VWcS7SqJCN3ApCqgbsVhal+F/Ps8qkaCcI6
zhb9hTKnhhF6+jIYou2l+zqSbUuA64eUz89myrSXfY2LxKRMWDa1NbSEwSifpehC
UwGaLcWvVO/cdMxR2k8RnrrXBse8G3AdQbPzjzKce2kIww+xvGZ4L5CaIRQFGZ28
Z00QJXN1kS+E32/zUjFZcgFqCVoq/pxk7yNv4yRGzNtIBoLRqZwrdA+xnInVz9Te
u1pr8GS+gdlrmyjblv9Nu61rBGO3P7ocfhDpvf1y6k49KI4ACEyd0UcXv28GIGL6
75NFRP23bCeSI0MowdtSGwDzk4fe6WsfN2IKbjODQad3E+ez4BRjiQKDfXdb/yPh
VWPXg8cV2docDVOJi/v29pwgzivYDTkkqJkx1PZjbt0/z97koIbhVhUI4xW4zclo
+v5st29W0IzkvLkGLl7Tk83B9G9GUdwpfzX4Ju+pFAQMhXr3UvoENno+EsUVSqqy
lSQE6eWejF+c8NBGSyP4bImiJTM+oofu5O/pzboZ1ADBSkTenubIEp7w1WMazBJO
L08YWXR89XjJLyWWsgKIjACidSsdElxFKPar8fv30W+j9iw87OQuE+apVryeH7g7
bik1gSL+0HVballIki8cODE1Ysm36yfDLWDQqgO0emC5GHPDbNiVyUhLLdSdUIqM
H6hpW7LH6PokcYAAYVmxja+ZZpsq9PDjejGrGI6FDtdrYHvH2qjC/IaFGpk21b2b
iet/YOscjRiGBC/g1I8KXrH05nIYeMNIJTRQxppz/wUv+sgs2Gxi6Fw9SoMZ34zv
5fyEDk2oLBFdZFzhb8KAupPYsWY+aQwcGu7FApyQvqqkZyz1CZ5jFzbJlkqOZ5Np
2Zdhf5x4xW5VENUY9antRgwfG/HsDgLXy/voN3Ir8swWUD/0prY7UZKbzb/sTsgq
BEsqVRQ2bqedgX6eQ7hsaZD85YkEh/9HKv2B9ZYBRQ5TyU7B2oeSMt/KniKfMFJW
RcQUmXD31GYouuZPg/lsOtsUQUX2j/oCWXAsfY2ZhAADQA7HtI+3lGL4pgW0h/e4
nJFW7wbhpYS5HbwfQxdQLRS6g7HMc86ef4MXTKG1URFNs3KWluWeZyXmJDEwdWxe
Ivs0eDB7wJZgBk7d48P0wiQ9geXs8WpfxMCw/ZssKyTUhs9VKXnf/Xzn6l+Opcfr
wxjemxitCf6pS/sPOthcE1CsY+YNo8ZNrwJJpf+mYQB9Ss0vA7UAqs5IMjjiANZ+
KtoICnaMTd4NJ+FrxMs7Ts7vzB5RS4CQz4SVeBNsBHmbLK6drg+YpUNmWsoQaWUt
7i6P1tTmVq0bjcnKDjez+TLxKNZoWdzDQZmGVpLBfQATkB1c6/lRs1A0VPAK6z+g
tFXadQPXjG5UJvf3TElNHHJYApfp0XtQ/YDgl4ebxBcKhiuUW4I2OsjSuxEp4v3v
DSbKqiGZEGegP72iLmmqZj6HR+VS6+XM1STXi+7WEFCuQpnLkcUlIvEh3jUlvHCX
K6wdfhoYW3ysLeHt3C+lf2C/u7Jq26ERyO9eP1G1Ot2kmdc3s1mfIGRGGblNwUtg
61lNP9TzEKrmFOfEq1rTbZWWmCM81IQV7ry/J7xHXB1zoxfzd69Mz94i/pm/ZsEQ
lWT/GFgrL/MeISIDGA8XtWL4y/kGiFHfW+W2XYP4f5SA2/LYt9bqWBpivPrKYxY5
2CKvIl2GTNR3qktAOwc1SqZ3e2PU5Jqn5qLhq+mwAuWWBySqC/rYBghISTNsFqnU
B/FFOuPNbWoc5QVNOkwwz0r5Z+ps6cHZoGIA2GUMzrl9zypo6wkWsIhmbJfKx4pM
jRl1puMzfyYWnZBLHEu9QZ2gEL4ci9ymXrZBQwQfhdlE/bTaRahklbt5R9UGylV5
XDcKMueZihujAivd6ECkdWAGzRHXzlbHUgD1cQJTS9yUA6Ud2xRLylKSBI/NvHQJ
8/a0zNydB/1KqrZJaU6S6R1pUH/BsAivCRjehuHwnMYiIh5QcybHOBA8058Wt1gs
Ur/Wqj8ffxMe48dfqU2dqKdCNI7oPHhM31gQtdUwMRQuidKcgpqtBF3VaBXXjBDx
P+TWY85+crgLeLRxm3DzZMR7h0CYPbb8pZgC61V0yOudAmtndSu/4ditqJ4hYVVK
nNIgus7tJanSMfkzYWDgQ5NY15glN+wRvX7EVwOSzzJb4/WO6zmmnb5AzoxrMyJs
F3OOo232GBf/dmIo0g/ODThhvr12Z831q40dnBTugZGS+CY1WfKrn+5y5Wg+0sDD
BwFT/P6tYs6UlsaW2VHKzRvdaNPJrfjqYDkoETmYjQ1I7yEBnbgjt+QBgJiCkhgW
KalLud9u09yrhElzqSz36tS2d7qP1OQtfMICebiMUp6mVZyMItGbdlOpRqwJfIM3
+XnGflJRydh4fL/4QVT8FkWxhylSUNOKlpsBhz70EjTPgq+Mh5v+FfjyCXYmh13y
gUwnYkd35SwZC0MHrewtT+fyWGPARpKoMuDk2abNAQkcfcieAzpsimjvmWDCrxe6
mXhT69T1TYKiFBIvuwDjZSinluROzcXMXSynzew5m5Zk7G3CZSRjiQ4i0/gr0UQ4
7VV9e9PGOgzM2V8MdfTcrZ2KTn01s8tAQD0oc264KE8dAqilqCTD2Q3x/T8L/1VU
XcfMoEm3cYedsTuKnjY4evL8LY9weyGbKMadfp6kAIlB+xE+dWiArd1N0/IVv+2u
oOrlWAd4slfP1paDj/TPzEa4KJVyP3ojxmhVRTjaKunf8ZFV0Np69S+KiWQND0D7
T5NMkObcjKJ/tcno4JWf/SeK4pCrWt9Czwv0PtomaMY=
`pragma protect end_protected
