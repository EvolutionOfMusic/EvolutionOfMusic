-- niosII_system.vhd

-- Generated using ACDS version 12.1sp1 243 at 2016.03.23.15:55:29

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosII_system is
	port (
		reset_0_reset_n                                  : in    std_logic                     := '0';             --                                     reset_0.reset_n
		spi_0_external_MISO                              : in    std_logic                     := '0';             --                              spi_0_external.MISO
		spi_0_external_MOSI                              : out   std_logic;                                        --                                            .MOSI
		spi_0_external_SCLK                              : out   std_logic;                                        --                                            .SCLK
		spi_0_external_SS_n                              : out   std_logic;                                        --                                            .SS_n
		up_clocks_0_sys_clk_reset_reset_n                : out   std_logic;                                        --                   up_clocks_0_sys_clk_reset.reset_n
		audio_0_external_interface_ADCDAT                : in    std_logic                     := '0';             --                  audio_0_external_interface.ADCDAT
		audio_0_external_interface_ADCLRCK               : in    std_logic                     := '0';             --                                            .ADCLRCK
		audio_0_external_interface_BCLK                  : in    std_logic                     := '0';             --                                            .BCLK
		audio_0_external_interface_DACDAT                : out   std_logic;                                        --                                            .DACDAT
		audio_0_external_interface_DACLRCK               : in    std_logic                     := '0';             --                                            .DACLRCK
		clk_1_clk_in_clk                                 : in    std_logic                     := '0';             --                                clk_1_clk_in.clk
		up_clocks_0_sdram_clk_clk                        : out   std_logic;                                        --                       up_clocks_0_sdram_clk.clk
		audio_and_video_config_0_external_interface_SDAT : inout std_logic                     := '0';             -- audio_and_video_config_0_external_interface.SDAT
		audio_and_video_config_0_external_interface_SCLK : out   std_logic;                                        --                                            .SCLK
		up_clocks_0_audio_clk_clk                        : out   std_logic;                                        --                       up_clocks_0_audio_clk.clk
		reset_reset_n                                    : in    std_logic                     := '0';             --                                       reset.reset_n
		sdram_0_wire_addr                                : out   std_logic_vector(11 downto 0);                    --                                sdram_0_wire.addr
		sdram_0_wire_ba                                  : out   std_logic_vector(1 downto 0);                     --                                            .ba
		sdram_0_wire_cas_n                               : out   std_logic;                                        --                                            .cas_n
		sdram_0_wire_cke                                 : out   std_logic;                                        --                                            .cke
		sdram_0_wire_cs_n                                : out   std_logic;                                        --                                            .cs_n
		sdram_0_wire_dq                                  : inout std_logic_vector(15 downto 0) := (others => '0'); --                                            .dq
		sdram_0_wire_dqm                                 : out   std_logic_vector(1 downto 0);                     --                                            .dqm
		sdram_0_wire_ras_n                               : out   std_logic;                                        --                                            .ras_n
		sdram_0_wire_we_n                                : out   std_logic;                                        --                                            .we_n
		clk_clk                                          : in    std_logic                     := '0';             --                                         clk.clk
		sram_0_external_interface_DQ                     : inout std_logic_vector(15 downto 0) := (others => '0'); --                   sram_0_external_interface.DQ
		sram_0_external_interface_ADDR                   : out   std_logic_vector(17 downto 0);                    --                                            .ADDR
		sram_0_external_interface_LB_N                   : out   std_logic;                                        --                                            .LB_N
		sram_0_external_interface_UB_N                   : out   std_logic;                                        --                                            .UB_N
		sram_0_external_interface_CE_N                   : out   std_logic;                                        --                                            .CE_N
		sram_0_external_interface_OE_N                   : out   std_logic;                                        --                                            .OE_N
		sram_0_external_interface_WE_N                   : out   std_logic                                         --                                            .WE_N
	);
end entity niosII_system;

architecture rtl of niosII_system is
	component niosII_system_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_begintransfer       : in  std_logic                     := 'X';             -- begintransfer
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_select              : in  std_logic                     := 'X';             -- chipselect
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component niosII_system_nios2_qsys_0;

	component niosII_system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			clken      : in  std_logic                     := 'X';             -- clken
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X'              -- reset
		);
	end component niosII_system_onchip_memory2_0;

	component niosII_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component niosII_system_sysid_qsys_0;

	component niosII_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component niosII_system_timer_0;

	component niosII_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component niosII_system_jtag_uart_0;

	component niosII_system_sdram_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component niosII_system_sdram_0;

	component niosII_system_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(17 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component niosII_system_sram_0;

	component niosII_system_gate_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component niosII_system_gate_timer;

	component niosII_system_audio_0 is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
			from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
			from_adc_left_channel_data   : out std_logic_vector(31 downto 0);                    -- data
			from_adc_left_channel_valid  : out std_logic;                                        -- valid
			from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
			from_adc_right_channel_data  : out std_logic_vector(31 downto 0);                    -- data
			from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_ADCDAT                   : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK                  : in  std_logic                     := 'X';             -- export
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component niosII_system_audio_0;

	component niosII_system_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component niosII_system_audio_and_video_config_0;

	component niosII_system_up_clocks_0 is
		port (
			CLOCK_50    : in  std_logic := 'X'; -- clk
			reset       : in  std_logic := 'X'; -- reset
			sys_clk     : out std_logic;        -- clk
			sys_reset_n : out std_logic;        -- reset_n
			SDRAM_CLK   : out std_logic;        -- clk
			CLOCK_27    : in  std_logic := 'X'; -- clk
			AUD_CLK     : out std_logic         -- clk
		);
	end component niosII_system_up_clocks_0;

	component niosII_system_synthesizer_0 is
		port (
			reset_n                    : in  std_logic                     := 'X';             -- reset_n
			avs_writedata_voice_select : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_write_n_voice_select   : in  std_logic                     := 'X';             -- write_n
			aso_ready_audio_in         : in  std_logic                     := 'X';             -- ready
			aso_data_audio_out         : out std_logic_vector(31 downto 0);                    -- data
			aso_valid_audio_out        : out std_logic;                                        -- valid
			csi_clk50M                 : in  std_logic                     := 'X';             -- clk
			csi_clk32k                 : in  std_logic                     := 'X'              -- clk
		);
	end component niosII_system_synthesizer_0;

	component niosII_system_spi_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component niosII_system_spi_0;

	component niosII_system_nios2_qsys_0_instruction_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component niosII_system_nios2_qsys_0_instruction_master_translator;

	component niosII_system_nios2_qsys_0_data_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_write          : in  std_logic                     := 'X';             -- write
			av_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess    : in  std_logic                     := 'X'              -- debugaccess
		);
	end component niosII_system_nios2_qsys_0_data_master_translator;

	component niosII_system_nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			av_address       : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_write         : in  std_logic                     := 'X';             -- write
			av_read          : in  std_logic                     := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest   : out std_logic;                                        -- waitrequest
			av_readdatavalid : out std_logic;                                        -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_lock          : in  std_logic                     := 'X';             -- lock
			cp_valid         : out std_logic;                                        -- valid
			cp_data          : out std_logic_vector(99 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                        -- startofpacket
			cp_endofpacket   : out std_logic;                                        -- endofpacket
			cp_ready         : in  std_logic                     := 'X';             -- ready
			rp_valid         : in  std_logic                     := 'X';             -- valid
			rp_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rp_ready         : out std_logic                                         -- ready
		);
	end component niosII_system_nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent;

	component niosII_system_nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			av_address       : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_write         : in  std_logic                     := 'X';             -- write
			av_read          : in  std_logic                     := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest   : out std_logic;                                        -- waitrequest
			av_readdatavalid : out std_logic;                                        -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_lock          : in  std_logic                     := 'X';             -- lock
			cp_valid         : out std_logic;                                        -- valid
			cp_data          : out std_logic_vector(99 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                        -- startofpacket
			cp_endofpacket   : out std_logic;                                        -- endofpacket
			cp_ready         : in  std_logic                     := 'X';             -- ready
			rp_valid         : in  std_logic                     := 'X';             -- valid
			rp_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rp_ready         : out std_logic                                         -- ready
		);
	end component niosII_system_nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent;

	component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(100 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component niosII_system_onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent;

	component niosII_system_sdram_0_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(81 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(82 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(15 downto 0)                     -- data
		);
	end component niosII_system_sdram_0_s1_translator_avalon_universal_slave_0_agent;

	component niosII_system_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(82 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component niosII_system_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component niosII_system_sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(81 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(82 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(15 downto 0)                     -- data
		);
	end component niosII_system_sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent;

	component niosII_system_sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(82 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component niosII_system_sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component niosII_system_audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent;

	component niosII_system_synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent;

	component niosII_system_spi_0_spi_control_port_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_spi_0_spi_control_port_translator_avalon_universal_slave_0_agent;

	component niosII_system_sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent;

	component niosII_system_timer_0_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_timer_0_s1_translator_avalon_universal_slave_0_agent;

	component niosII_system_jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent;

	component niosII_system_gate_timer_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                      -- data
		);
	end component niosII_system_gate_timer_s1_translator_avalon_universal_slave_0_agent;

	component niosII_system_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component niosII_system_addr_router;

	component niosII_system_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component niosII_system_addr_router_001;

	component niosII_system_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component niosII_system_id_router;

	component niosII_system_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(81 downto 0);                    -- data
			src_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component niosII_system_id_router_002;

	component niosII_system_id_router_007 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component niosII_system_id_router_007;

	component niosII_system_burst_adapter is
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(81 downto 0);                    -- data
			source0_channel       : out std_logic_vector(10 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component niosII_system_burst_adapter;

	component niosII_system_rst_controller is
		port (
			reset_in0 : in  std_logic := 'X'; -- reset
			reset_in1 : in  std_logic := 'X'; -- reset
			clk       : in  std_logic := 'X'; -- clk
			reset_out : out std_logic         -- reset
		);
	end component niosII_system_rst_controller;

	component niosII_system_rst_controller_001 is
		port (
			reset_in0 : in  std_logic := 'X'; -- reset
			clk       : in  std_logic := 'X'; -- clk
			reset_out : out std_logic         -- reset
		);
	end component niosII_system_rst_controller_001;

	component niosII_system_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(99 downto 0);                    -- data
			src2_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(99 downto 0);                    -- data
			src3_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(99 downto 0);                    -- data
			src4_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic;                                        -- endofpacket
			src5_ready         : in  std_logic                     := 'X';             -- ready
			src5_valid         : out std_logic;                                        -- valid
			src5_data          : out std_logic_vector(99 downto 0);                    -- data
			src5_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src5_startofpacket : out std_logic;                                        -- startofpacket
			src5_endofpacket   : out std_logic;                                        -- endofpacket
			src6_ready         : in  std_logic                     := 'X';             -- ready
			src6_valid         : out std_logic;                                        -- valid
			src6_data          : out std_logic_vector(99 downto 0);                    -- data
			src6_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src6_startofpacket : out std_logic;                                        -- startofpacket
			src6_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component niosII_system_cmd_xbar_demux;

	component niosII_system_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(99 downto 0);                    -- data
			src0_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(99 downto 0);                    -- data
			src1_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(99 downto 0);                    -- data
			src2_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(99 downto 0);                    -- data
			src3_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(99 downto 0);                    -- data
			src4_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(99 downto 0);                    -- data
			src5_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(99 downto 0);                    -- data
			src6_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(99 downto 0);                    -- data
			src7_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(99 downto 0);                    -- data
			src8_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(99 downto 0);                    -- data
			src9_channel        : out std_logic_vector(10 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(99 downto 0);                    -- data
			src10_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component niosII_system_cmd_xbar_demux_001;

	component niosII_system_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component niosII_system_cmd_xbar_mux;

	component niosII_system_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component niosII_system_rsp_xbar_demux;

	component niosII_system_rsp_xbar_demux_007 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(10 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component niosII_system_rsp_xbar_demux_007;

	component niosII_system_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                        -- ready
			sink5_valid         : in  std_logic                     := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                        -- ready
			sink6_valid         : in  std_logic                     := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component niosII_system_rsp_xbar_mux;

	component niosII_system_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(99 downto 0);                    -- data
			src_channel          : out std_logic_vector(10 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component niosII_system_rsp_xbar_mux_001;

	component niosII_system_width_adapter is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_ready          : out std_logic;                                        -- ready
			in_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			out_endofpacket   : out std_logic;                                        -- endofpacket
			out_data          : out std_logic_vector(81 downto 0);                    -- data
			out_channel       : out std_logic_vector(10 downto 0);                    -- channel
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic                                         -- startofpacket
		);
	end component niosII_system_width_adapter;

	component niosII_system_width_adapter_001 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_channel        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- channel
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_ready          : out std_logic;                                        -- ready
			in_data           : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			out_endofpacket   : out std_logic;                                        -- endofpacket
			out_data          : out std_logic_vector(99 downto 0);                    -- data
			out_channel       : out std_logic_vector(10 downto 0);                    -- channel
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic                                         -- startofpacket
		);
	end component niosII_system_width_adapter_001;

	component niosII_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component niosII_system_irq_mapper;

	component niosii_system_nios2_qsys_0_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(8 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect         : out std_logic;                                        -- chipselect
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_read               : out std_logic;                                        -- read
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_nios2_qsys_0_jtag_debug_module_translator;

	component niosii_system_onchip_memory2_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(11 downto 0);                    -- address
			av_write              : out std_logic;                                        -- write
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			av_read               : out std_logic;                                        -- read
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_onchip_memory2_0_s1_translator;

	component niosii_system_sdram_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(21 downto 0);                    -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable         : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect         : out std_logic;                                        -- chipselect
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable    : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_sdram_0_s1_translator;

	component niosii_system_sram_0_avalon_sram_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(17 downto 0);                    -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable         : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_sram_0_avalon_sram_slave_translator;

	component niosii_system_audio_and_video_config_0_avalon_av_config_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(1 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_audio_and_video_config_0_avalon_av_config_slave_translator;

	component niosii_system_synthesizer_0_voice_select_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_write              : out std_logic;                                        -- write
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_address            : out std_logic_vector(0 downto 0);                     -- address
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_chipselect         : out std_logic;                                        -- chipselect
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_synthesizer_0_voice_select_translator;

	component niosii_system_spi_0_spi_control_port_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(2 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect         : out std_logic;                                        -- chipselect
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_spi_0_spi_control_port_translator;

	component niosii_system_timer_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(2 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_readdata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect         : out std_logic;                                        -- chipselect
			av_read               : out std_logic;                                        -- read
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable    : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_timer_0_s1_translator;

	component niosii_system_jtag_uart_0_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			uav_address           : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read              : in  std_logic                     := 'X';             -- read
			uav_write             : in  std_logic                     := 'X';             -- write
			uav_waitrequest       : out std_logic;                                        -- waitrequest
			uav_readdatavalid     : out std_logic;                                        -- readdatavalid
			uav_byteenable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock              : in  std_logic                     := 'X';             -- lock
			uav_debugaccess       : in  std_logic                     := 'X';             -- debugaccess
			av_address            : out std_logic_vector(0 downto 0);                     -- address
			av_write              : out std_logic;                                        -- write
			av_read               : out std_logic;                                        -- read
			av_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect         : out std_logic;                                        -- chipselect
			av_begintransfer      : out std_logic;                                        -- begintransfer
			av_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			av_burstcount         : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable         : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable    : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock               : out std_logic;                                        -- lock
			av_clken              : out std_logic;                                        -- clken
			uav_clken             : in  std_logic                     := 'X';             -- clken
			av_debugaccess        : out std_logic;                                        -- debugaccess
			av_outputenable       : out std_logic                                         -- outputenable
		);
	end component niosii_system_jtag_uart_0_avalon_jtag_slave_translator;

	signal nios2_qsys_0_jtag_debug_module_reset_reset                                                                           : std_logic;                      -- nios2_qsys_0:jtag_debug_module_resetrequest -> [audio_and_video_config_0:reset, audio_and_video_config_0_avalon_av_config_slave_translator:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, nios2_qsys_0_jtag_debug_module_reset_reset:in, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rst_controller:reset_in1, rst_controller_002:reset_in0, spi_0_spi_control_port_translator:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, synthesizer_0_voice_select_translator:reset, synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:reset, synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal up_clocks_0_sys_clk_clk                                                                                              : std_logic;                      -- up_clocks_0:sys_clk -> [addr_router:clk, addr_router_001:clk, audio_0:clk, audio_and_video_config_0:clk, audio_and_video_config_0_avalon_av_config_slave_translator:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_004:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_006:clk, gate_timer:clk, gate_timer_s1_translator:clk, gate_timer_s1_translator_avalon_universal_slave_0_agent:clk, gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, rst_controller_001:clk, sdram_0:clk, sdram_0_s1_translator:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, spi_0:clk, spi_0_spi_control_port_translator:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sram_0:clk, sram_0_avalon_sram_slave_translator:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, synthesizer_0:csi_clk32k, synthesizer_0:csi_clk50M, synthesizer_0_voice_select_translator:clk, synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:clk, synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys_0:clock, sysid_qsys_0_control_slave_translator:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk]
	signal synthesizer_0_audio_valid                                                                                            : std_logic;                      -- synthesizer_0:aso_valid_audio_out -> audio_0:to_dac_left_channel_valid
	signal synthesizer_0_audio_data                                                                                             : std_logic_vector(31 downto 0);  -- synthesizer_0:aso_data_audio_out -> audio_0:to_dac_left_channel_data
	signal synthesizer_0_audio_ready                                                                                            : std_logic;                      -- audio_0:to_dac_left_channel_ready -> synthesizer_0:aso_ready_audio_in
	signal nios2_qsys_0_instruction_master_waitrequest                                                                          : std_logic;                      -- nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                                                                              : std_logic_vector(24 downto 0);  -- nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	signal nios2_qsys_0_instruction_master_read                                                                                 : std_logic;                      -- nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	signal nios2_qsys_0_instruction_master_readdata                                                                             : std_logic_vector(31 downto 0);  -- nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_data_master_waitrequest                                                                                 : std_logic;                      -- nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_writedata                                                                                   : std_logic_vector(31 downto 0);  -- nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	signal nios2_qsys_0_data_master_address                                                                                     : std_logic_vector(24 downto 0);  -- nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	signal nios2_qsys_0_data_master_write                                                                                       : std_logic;                      -- nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	signal nios2_qsys_0_data_master_read                                                                                        : std_logic;                      -- nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	signal nios2_qsys_0_data_master_readdata                                                                                    : std_logic_vector(31 downto 0);  -- nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_debugaccess                                                                                 : std_logic;                      -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	signal nios2_qsys_0_data_master_byteenable                                                                                  : std_logic_vector(3 downto 0);   -- nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(31 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address                                                : std_logic_vector(8 downto 0);   -- nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator:av_chipselect -> nios2_qsys_0:jtag_debug_module_select
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write                                                  : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0);  -- nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer                                          : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator:av_begintransfer -> nios2_qsys_0:jtag_debug_module_begintransfer
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                            : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                             : std_logic_vector(3 downto 0);   -- nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata                                                         : std_logic_vector(31 downto 0);  -- onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_address                                                           : std_logic_vector(11 downto 0);  -- onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect                                                        : std_logic;                      -- onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken                                                             : std_logic;                      -- onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_write                                                             : std_logic;                      -- onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata                                                          : std_logic_vector(31 downto 0);  -- onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable                                                        : std_logic_vector(3 downto 0);   -- onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	signal sdram_0_s1_translator_avalon_anti_slave_0_waitrequest                                                                : std_logic;                      -- sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	signal sdram_0_s1_translator_avalon_anti_slave_0_writedata                                                                  : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	signal sdram_0_s1_translator_avalon_anti_slave_0_address                                                                    : std_logic_vector(21 downto 0);  -- sdram_0_s1_translator:av_address -> sdram_0:az_addr
	signal sdram_0_s1_translator_avalon_anti_slave_0_chipselect                                                                 : std_logic;                      -- sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	signal sdram_0_s1_translator_avalon_anti_slave_0_write                                                                      : std_logic;                      -- sdram_0_s1_translator:av_write -> sdram_0_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_0_s1_translator_avalon_anti_slave_0_read                                                                       : std_logic;                      -- sdram_0_s1_translator:av_read -> sdram_0_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_0_s1_translator_avalon_anti_slave_0_readdata                                                                   : std_logic_vector(15 downto 0);  -- sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	signal sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid                                                              : std_logic;                      -- sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	signal sdram_0_s1_translator_avalon_anti_slave_0_byteenable                                                                 : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator:av_byteenable -> sdram_0_s1_translator_avalon_anti_slave_0_byteenable:in
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(15 downto 0);  -- sram_0_avalon_sram_slave_translator:av_writedata -> sram_0:writedata
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(17 downto 0);  -- sram_0_avalon_sram_slave_translator:av_address -> sram_0:address
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- sram_0_avalon_sram_slave_translator:av_write -> sram_0:write
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read                                                         : std_logic;                      -- sram_0_avalon_sram_slave_translator:av_read -> sram_0:read
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(15 downto 0);  -- sram_0:readdata -> sram_0_avalon_sram_slave_translator:av_readdata
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid                                                : std_logic;                      -- sram_0:readdatavalid -> sram_0_avalon_sram_slave_translator:av_readdatavalid
	signal sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable                                                   : std_logic_vector(1 downto 0);   -- sram_0_avalon_sram_slave_translator:av_byteenable -> sram_0:byteenable
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- audio_and_video_config_0:waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator:av_waitrequest
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- audio_and_video_config_0_avalon_av_config_slave_translator:av_writedata -> audio_and_video_config_0:writedata
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(1 downto 0);   -- audio_and_video_config_0_avalon_av_config_slave_translator:av_address -> audio_and_video_config_0:address
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator:av_write -> audio_and_video_config_0:write
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator:av_read -> audio_and_video_config_0:read
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- audio_and_video_config_0:readdata -> audio_and_video_config_0_avalon_av_config_slave_translator:av_readdata
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- audio_and_video_config_0_avalon_av_config_slave_translator:av_byteenable -> audio_and_video_config_0:byteenable
	signal synthesizer_0_voice_select_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0);  -- synthesizer_0_voice_select_translator:av_writedata -> synthesizer_0:avs_writedata_voice_select
	signal synthesizer_0_voice_select_translator_avalon_anti_slave_0_write                                                      : std_logic;                      -- synthesizer_0_voice_select_translator:av_write -> synthesizer_0_voice_select_translator_avalon_anti_slave_0_write:in
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata                                                      : std_logic_vector(31 downto 0);  -- spi_0_spi_control_port_translator:av_writedata -> spi_0:data_from_cpu
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_address                                                        : std_logic_vector(2 downto 0);   -- spi_0_spi_control_port_translator:av_address -> spi_0:mem_addr
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect                                                     : std_logic;                      -- spi_0_spi_control_port_translator:av_chipselect -> spi_0:spi_select
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_write                                                          : std_logic;                      -- spi_0_spi_control_port_translator:av_write -> spi_0_spi_control_port_translator_avalon_anti_slave_0_write:in
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_read                                                           : std_logic;                      -- spi_0_spi_control_port_translator:av_read -> spi_0_spi_control_port_translator_avalon_anti_slave_0_read:in
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata                                                       : std_logic_vector(31 downto 0);  -- spi_0:data_to_cpu -> spi_0_spi_control_port_translator:av_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(0 downto 0);   -- sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0);  -- sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                                                  : std_logic_vector(15 downto 0);  -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                                                    : std_logic_vector(2 downto 0);   -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                                                 : std_logic;                      -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                                                      : std_logic;                      -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                                                   : std_logic_vector(15 downto 0);  -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                             : std_logic;                      -- jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(0 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                                   : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                                    : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	signal gate_timer_s1_translator_avalon_anti_slave_0_writedata                                                               : std_logic_vector(15 downto 0);  -- gate_timer_s1_translator:av_writedata -> gate_timer:writedata
	signal gate_timer_s1_translator_avalon_anti_slave_0_address                                                                 : std_logic_vector(2 downto 0);   -- gate_timer_s1_translator:av_address -> gate_timer:address
	signal gate_timer_s1_translator_avalon_anti_slave_0_chipselect                                                              : std_logic;                      -- gate_timer_s1_translator:av_chipselect -> gate_timer:chipselect
	signal gate_timer_s1_translator_avalon_anti_slave_0_write                                                                   : std_logic;                      -- gate_timer_s1_translator:av_write -> gate_timer_s1_translator_avalon_anti_slave_0_write:in
	signal gate_timer_s1_translator_avalon_anti_slave_0_readdata                                                                : std_logic_vector(15 downto 0);  -- gate_timer:readdata -> gate_timer_s1_translator:av_readdata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest                                     : std_logic;                      -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount                                      : std_logic_vector(2 downto 0);   -- nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata                                       : std_logic_vector(31 downto 0);  -- nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address                                         : std_logic_vector(24 downto 0);  -- nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock                                            : std_logic;                      -- nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write                                           : std_logic;                      -- nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read                                            : std_logic;                      -- nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata                                        : std_logic_vector(31 downto 0);  -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess                                     : std_logic;                      -- nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable                                      : std_logic_vector(3 downto 0);   -- nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid                                   : std_logic;                      -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest                                            : std_logic;                      -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount                                             : std_logic_vector(2 downto 0);   -- nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata                                              : std_logic_vector(31 downto 0);  -- nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_address                                                : std_logic_vector(24 downto 0);  -- nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock                                                   : std_logic;                      -- nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_write                                                  : std_logic;                      -- nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_read                                                   : std_logic;                      -- nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata                                               : std_logic_vector(31 downto 0);  -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess                                            : std_logic;                      -- nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable                                             : std_logic_vector(3 downto 0);   -- nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid                                          : std_logic;                      -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);   -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(24 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);   -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(100 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(100 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(31 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                         : std_logic;                      -- onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                          : std_logic_vector(2 downto 0);   -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                           : std_logic_vector(31 downto 0);  -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                             : std_logic_vector(24 downto 0);  -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                               : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                            : std_logic_vector(31 downto 0);  -- onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                       : std_logic;                      -- onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                         : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                          : std_logic_vector(3 downto 0);   -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                  : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                        : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                         : std_logic_vector(100 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                        : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                               : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                     : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                             : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                      : std_logic_vector(100 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                     : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                   : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                    : std_logic_vector(31 downto 0);  -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                   : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                  : std_logic;                      -- sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                   : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                    : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                                      : std_logic_vector(24 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                                        : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                         : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                         : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                     : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                : std_logic;                      -- sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                  : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                   : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                           : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                 : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                         : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                  : std_logic_vector(82 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                 : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                        : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                              : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                      : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                               : std_logic_vector(82 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                              : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                            : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                             : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                            : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- sram_0_avalon_sram_slave_translator:uav_waitrequest -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(1 downto 0);   -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_sram_slave_translator:uav_burstcount
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(15 downto 0);  -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_sram_slave_translator:uav_writedata
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_sram_slave_translator:uav_address
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_sram_slave_translator:uav_write
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_sram_slave_translator:uav_lock
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_sram_slave_translator:uav_read
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(15 downto 0);  -- sram_0_avalon_sram_slave_translator:uav_readdata -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- sram_0_avalon_sram_slave_translator:uav_readdatavalid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_sram_slave_translator:uav_debugaccess
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(1 downto 0);   -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_sram_slave_translator:uav_byteenable
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(82 downto 0);  -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(82 downto 0);  -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(15 downto 0);  -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator:uav_waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_burstcount
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_writedata
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(24 downto 0);  -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_address
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_write
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_lock
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_read
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdata -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdatavalid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_debugaccess
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_byteenable
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(100 downto 0); -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(100 downto 0); -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(31 downto 0);  -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- synthesizer_0_voice_select_translator:uav_waitrequest -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);   -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_burstcount -> synthesizer_0_voice_select_translator:uav_burstcount
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0);  -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_writedata -> synthesizer_0_voice_select_translator:uav_writedata
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(24 downto 0);  -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_address -> synthesizer_0_voice_select_translator:uav_address
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_write -> synthesizer_0_voice_select_translator:uav_write
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_lock -> synthesizer_0_voice_select_translator:uav_lock
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_read -> synthesizer_0_voice_select_translator:uav_read
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0);  -- synthesizer_0_voice_select_translator:uav_readdata -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_readdata
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- synthesizer_0_voice_select_translator:uav_readdatavalid -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_debugaccess -> synthesizer_0_voice_select_translator:uav_debugaccess
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);   -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:m0_byteenable -> synthesizer_0_voice_select_translator:uav_byteenable
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_source_valid -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(100 downto 0); -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_source_data -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(100 downto 0); -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rf_sink_ready -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(31 downto 0);  -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest                                      : std_logic;                      -- spi_0_spi_control_port_translator:uav_waitrequest -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount                                       : std_logic_vector(2 downto 0);   -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_0_spi_control_port_translator:uav_burstcount
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata                                        : std_logic_vector(31 downto 0);  -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_0_spi_control_port_translator:uav_writedata
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address                                          : std_logic_vector(24 downto 0);  -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> spi_0_spi_control_port_translator:uav_address
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write                                            : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> spi_0_spi_control_port_translator:uav_write
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock                                             : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> spi_0_spi_control_port_translator:uav_lock
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read                                             : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> spi_0_spi_control_port_translator:uav_read
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata                                         : std_logic_vector(31 downto 0);  -- spi_0_spi_control_port_translator:uav_readdata -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                    : std_logic;                      -- spi_0_spi_control_port_translator:uav_readdatavalid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess                                      : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_0_spi_control_port_translator:uav_debugaccess
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable                                       : std_logic_vector(3 downto 0);   -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_0_spi_control_port_translator:uav_byteenable
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                               : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid                                     : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                             : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data                                      : std_logic_vector(100 downto 0); -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready                                     : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                            : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                  : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                          : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                   : std_logic_vector(100 downto 0); -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                  : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                 : std_logic_vector(31 downto 0);  -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);   -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(24 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);   -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(100 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(100 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                  : std_logic;                      -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                   : std_logic_vector(2 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                    : std_logic_vector(31 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                                      : std_logic_vector(24 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                         : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                         : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                     : std_logic_vector(31 downto 0);  -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                : std_logic;                      -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                  : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                   : std_logic_vector(3 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                           : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                 : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                         : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                  : std_logic_vector(100 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                 : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                      : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                               : std_logic_vector(100 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                            : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                             : std_logic_vector(31 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                            : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(24 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(100 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(100 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                               : std_logic;                      -- gate_timer_s1_translator:uav_waitrequest -> gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                : std_logic_vector(2 downto 0);   -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> gate_timer_s1_translator:uav_burstcount
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                 : std_logic_vector(31 downto 0);  -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> gate_timer_s1_translator:uav_writedata
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_address                                                   : std_logic_vector(24 downto 0);  -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> gate_timer_s1_translator:uav_address
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_write                                                     : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> gate_timer_s1_translator:uav_write
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                      : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> gate_timer_s1_translator:uav_lock
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_read                                                      : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> gate_timer_s1_translator:uav_read
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                  : std_logic_vector(31 downto 0);  -- gate_timer_s1_translator:uav_readdata -> gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                             : std_logic;                      -- gate_timer_s1_translator:uav_readdatavalid -> gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                               : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> gate_timer_s1_translator:uav_debugaccess
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                : std_logic_vector(3 downto 0);   -- gate_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> gate_timer_s1_translator:uav_byteenable
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                        : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                              : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                      : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                               : std_logic_vector(100 downto 0); -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                              : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                     : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                           : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                   : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                            : std_logic_vector(100 downto 0); -- gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                           : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                         : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                          : std_logic_vector(31 downto 0);  -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                         : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                            : std_logic;                      -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                                  : std_logic;                      -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                          : std_logic;                      -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data                                   : std_logic_vector(99 downto 0);  -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                                  : std_logic;                      -- addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                   : std_logic;                      -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid                                         : std_logic;                      -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                 : std_logic;                      -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data                                          : std_logic_vector(99 downto 0);  -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready                                         : std_logic;                      -- addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(99 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                      -- id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                         : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                               : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                       : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                : std_logic_vector(99 downto 0);  -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                               : std_logic;                      -- id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                  : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                        : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                         : std_logic_vector(81 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                        : std_logic;                      -- id_router_002:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(81 downto 0);  -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_003:sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(99 downto 0);  -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_004:sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(99 downto 0);  -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_005:sink_ready -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:rp_ready
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket                                      : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid                                            : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket                                    : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data                                             : std_logic_vector(99 downto 0);  -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready                                            : std_logic;                      -- id_router_006:sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(99 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_007:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                  : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                         : std_logic_vector(99 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                        : std_logic;                      -- id_router_008:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(99 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                      -- id_router_009:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                               : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                     : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                             : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_data                                                      : std_logic_vector(99 downto 0);  -- gate_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                     : std_logic;                      -- id_router_010:sink_ready -> gate_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal burst_adapter_source0_endofpacket                                                                                    : std_logic;                      -- burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                                          : std_logic;                      -- burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                                  : std_logic;                      -- burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                                           : std_logic_vector(81 downto 0);  -- burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                                          : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                                        : std_logic_vector(10 downto 0);  -- burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                                                : std_logic;                      -- burst_adapter_001:source0_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                                      : std_logic;                      -- burst_adapter_001:source0_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                                              : std_logic;                      -- burst_adapter_001:source0_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                                       : std_logic_vector(81 downto 0);  -- burst_adapter_001:source0_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                                      : std_logic;                      -- sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                                    : std_logic_vector(10 downto 0);  -- burst_adapter_001:source0_channel -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                                       : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, gate_timer_s1_translator:reset, gate_timer_s1_translator_avalon_universal_slave_0_agent:reset, gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, irq_mapper:reset, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram_0:reset, sram_0_avalon_sram_slave_translator:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	signal rst_controller_001_reset_out_reset                                                                                   : std_logic;                      -- rst_controller_001:reset_out -> audio_0:reset
	signal rst_controller_002_reset_out_reset                                                                                   : std_logic;                      -- rst_controller_002:reset_out -> up_clocks_0:reset
	signal cmd_xbar_demux_src0_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                                            : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                                            : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                                            : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_src3_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                                            : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_src4_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_src4_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_src4_ready                                                                                            : std_logic;                      -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	signal cmd_xbar_demux_src5_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	signal cmd_xbar_demux_src5_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	signal cmd_xbar_demux_src5_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	signal cmd_xbar_demux_src5_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	signal cmd_xbar_demux_src5_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	signal cmd_xbar_demux_src5_ready                                                                                            : std_logic;                      -- cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	signal cmd_xbar_demux_src6_endofpacket                                                                                      : std_logic;                      -- cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	signal cmd_xbar_demux_src6_valid                                                                                            : std_logic;                      -- cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	signal cmd_xbar_demux_src6_startofpacket                                                                                    : std_logic;                      -- cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	signal cmd_xbar_demux_src6_data                                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	signal cmd_xbar_demux_src6_channel                                                                                          : std_logic_vector(10 downto 0);  -- cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	signal cmd_xbar_demux_src6_ready                                                                                            : std_logic;                      -- cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                                        : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_001_src4_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_001_src4_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	signal cmd_xbar_demux_001_src5_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	signal cmd_xbar_demux_001_src5_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	signal cmd_xbar_demux_001_src5_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	signal cmd_xbar_demux_001_src6_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	signal cmd_xbar_demux_001_src6_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	signal cmd_xbar_demux_001_src6_ready                                                                                        : std_logic;                      -- cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	signal cmd_xbar_demux_001_src7_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src7_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src7_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src8_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src8_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src8_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src8_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src8_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                                                  : std_logic;                      -- cmd_xbar_demux_001:src9_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src9_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_001:src9_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                                         : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src9_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                                      : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src9_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src10_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src10_endofpacket -> gate_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_001:src10_valid -> gate_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_001:src10_startofpacket -> gate_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                                        : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src10_data -> gate_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src10_channel                                                                                     : std_logic_vector(10 downto 0);  -- cmd_xbar_demux_001:src10_channel -> gate_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                                      : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                                            : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                                    : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                                             : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                                          : std_logic_vector(10 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                                            : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                                      : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                                            : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                                    : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                                             : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                                          : std_logic_vector(10 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                                            : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_005_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_006_src1_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src1_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src1_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src1_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src1_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src1_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                                  : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                                        : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                                : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                                         : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                                      : std_logic_vector(10 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal addr_router_src_endofpacket                                                                                          : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                                : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                                        : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                                 : std_logic_vector(99 downto 0);  -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                              : std_logic_vector(10 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                                : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                                         : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                               : std_logic;                      -- rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                                       : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                                : std_logic_vector(99 downto 0);  -- rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                                             : std_logic_vector(10 downto 0);  -- rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                               : std_logic;                      -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                                      : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                                            : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                                    : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                                             : std_logic_vector(99 downto 0);  -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                                          : std_logic_vector(10 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                                            : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                                     : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                                           : std_logic;                      -- rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                                   : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                                            : std_logic_vector(99 downto 0);  -- rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                                           : std_logic;                      -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                                         : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                               : std_logic;                      -- cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                                       : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                                : std_logic_vector(99 downto 0);  -- cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                                             : std_logic_vector(10 downto 0);  -- cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                               : std_logic;                      -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                                            : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                                  : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                                          : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                                   : std_logic_vector(99 downto 0);  -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                                : std_logic_vector(10 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                                  : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                                           : std_logic;                      -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                                        : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                                              : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                                      : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux_004:src_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux_004:src_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux_004:src_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_004:src_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- cmd_xbar_mux_004:src_channel -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                                           : std_logic;                      -- audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                                        : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                              : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                                      : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_mux_005_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux_005:src_endofpacket -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_005_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux_005:src_valid -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_005_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux_005:src_startofpacket -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_005_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_005:src_data -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_005_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- cmd_xbar_mux_005:src_channel -> synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_005_src_ready                                                                                           : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	signal id_router_005_src_endofpacket                                                                                        : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                              : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                                      : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_mux_006_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux_006:src_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_006_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux_006:src_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_006_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux_006:src_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_006_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_006:src_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_006_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- cmd_xbar_mux_006:src_channel -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_006_src_ready                                                                                           : std_logic;                      -- spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	signal id_router_006_src_endofpacket                                                                                        : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                              : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                                      : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                                        : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                                        : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                              : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                                      : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                                        : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                              : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                                      : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                                        : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                              : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                                      : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_001_src10_ready                                                                                       : std_logic;                      -- gate_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	signal id_router_010_src_endofpacket                                                                                        : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                                              : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                                      : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                               : std_logic_vector(99 downto 0);  -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                                              : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_002:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_002_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_002_src_ready                                                                                           : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	signal width_adapter_src_endofpacket                                                                                        : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                                              : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                                      : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                                               : std_logic_vector(81 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                                              : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_002_src_endofpacket                                                                                        : std_logic;                      -- id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_002_src_valid                                                                                              : std_logic;                      -- id_router_002:src_valid -> width_adapter_001:in_valid
	signal id_router_002_src_startofpacket                                                                                      : std_logic;                      -- id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_002_src_data                                                                                               : std_logic_vector(81 downto 0);  -- id_router_002:src_data -> width_adapter_001:in_data
	signal id_router_002_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_002:src_channel -> width_adapter_001:in_channel
	signal id_router_002_src_ready                                                                                              : std_logic;                      -- width_adapter_001:in_ready -> id_router_002:src_ready
	signal width_adapter_001_src_endofpacket                                                                                    : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal width_adapter_001_src_valid                                                                                          : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	signal width_adapter_001_src_startofpacket                                                                                  : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal width_adapter_001_src_data                                                                                           : std_logic_vector(99 downto 0);  -- width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	signal width_adapter_001_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                                        : std_logic_vector(10 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	signal cmd_xbar_mux_003_src_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                                           : std_logic;                      -- cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                                            : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	signal cmd_xbar_mux_003_src_channel                                                                                         : std_logic_vector(10 downto 0);  -- cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	signal cmd_xbar_mux_003_src_ready                                                                                           : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	signal width_adapter_002_src_endofpacket                                                                                    : std_logic;                      -- width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal width_adapter_002_src_valid                                                                                          : std_logic;                      -- width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	signal width_adapter_002_src_startofpacket                                                                                  : std_logic;                      -- width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal width_adapter_002_src_data                                                                                           : std_logic_vector(81 downto 0);  -- width_adapter_002:out_data -> burst_adapter_001:sink0_data
	signal width_adapter_002_src_ready                                                                                          : std_logic;                      -- burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                                        : std_logic_vector(10 downto 0);  -- width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	signal id_router_003_src_endofpacket                                                                                        : std_logic;                      -- id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	signal id_router_003_src_valid                                                                                              : std_logic;                      -- id_router_003:src_valid -> width_adapter_003:in_valid
	signal id_router_003_src_startofpacket                                                                                      : std_logic;                      -- id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	signal id_router_003_src_data                                                                                               : std_logic_vector(81 downto 0);  -- id_router_003:src_data -> width_adapter_003:in_data
	signal id_router_003_src_channel                                                                                            : std_logic_vector(10 downto 0);  -- id_router_003:src_channel -> width_adapter_003:in_channel
	signal id_router_003_src_ready                                                                                              : std_logic;                      -- width_adapter_003:in_ready -> id_router_003:src_ready
	signal width_adapter_003_src_endofpacket                                                                                    : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal width_adapter_003_src_valid                                                                                          : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	signal width_adapter_003_src_startofpacket                                                                                  : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal width_adapter_003_src_data                                                                                           : std_logic_vector(99 downto 0);  -- width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	signal width_adapter_003_src_ready                                                                                          : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                                        : std_logic_vector(10 downto 0);  -- width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	signal irq_mapper_receiver0_irq                                                                                             : std_logic;                      -- timer_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                                             : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                                             : std_logic;                      -- gate_timer:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                                             : std_logic;                      -- spi_0:irq -> irq_mapper:receiver3_irq
	signal nios2_qsys_0_d_irq_irq                                                                                               : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal reset_reset_n_ports_inv                                                                                              : std_logic;                      -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal nios2_qsys_0_jtag_debug_module_reset_reset_ports_inv                                                                 : std_logic;                      -- nios2_qsys_0_jtag_debug_module_reset_reset:inv -> [spi_0:reset_n, synthesizer_0:reset_n]
	signal sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                                            : std_logic;                      -- sdram_0_s1_translator_avalon_anti_slave_0_write:inv -> sdram_0:az_wr_n
	signal sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv                                                             : std_logic;                      -- sdram_0_s1_translator_avalon_anti_slave_0_read:inv -> sdram_0:az_rd_n
	signal sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                                       : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram_0:az_be_n
	signal synthesizer_0_voice_select_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                      -- synthesizer_0_voice_select_translator_avalon_anti_slave_0_write:inv -> synthesizer_0:avs_write_n_voice_select
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv                                                : std_logic;                      -- spi_0_spi_control_port_translator_avalon_anti_slave_0_write:inv -> spi_0:write_n
	signal spi_0_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv                                                 : std_logic;                      -- spi_0_spi_control_port_translator_avalon_anti_slave_0_read:inv -> spi_0:read_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                                            : std_logic;                      -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_0:av_write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                                          : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_0:av_read_n
	signal gate_timer_s1_translator_avalon_anti_slave_0_write_ports_inv                                                         : std_logic;                      -- gate_timer_s1_translator_avalon_anti_slave_0_write:inv -> gate_timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                                             : std_logic;                      -- rst_controller_reset_out_reset:inv -> [gate_timer:reset_n, jtag_uart_0:rst_n, nios2_qsys_0:reset_n, sdram_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]

begin

	nios2_qsys_0 : component niosII_system_nios2_qsys_0
		port map (
			clk                                   => up_clocks_0_sys_clk_clk,                                                     --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                    --                   reset_n.reset_n
			d_address                             => nios2_qsys_0_data_master_address,                                            --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                                         --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                               --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                                           --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                                        --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                                              --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                                          --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                                        --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                                     --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                                        --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                                    --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                                 --                          .waitrequest
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                                      --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                                  --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address,       --         jtag_debug_module.address
			jtag_debug_module_begintransfer       => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer, --                          .begintransfer
			jtag_debug_module_byteenable          => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,    --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,   --                          .debugaccess
			jtag_debug_module_readdata            => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,      --                          .readdata
			jtag_debug_module_select              => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect,    --                          .chipselect
			jtag_debug_module_write               => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write,         --                          .write
			jtag_debug_module_writedata           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,     --                          .writedata
			no_ci_readra                          => open                                                                         -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component niosII_system_onchip_memory2_0
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                       --   clk1.clk
			address    => onchip_memory2_0_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			chipselect => onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			clken      => onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			readdata   => onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			write      => onchip_memory2_0_s1_translator_avalon_anti_slave_0_write,      --       .write
			writedata  => onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset                                 -- reset1.reset
		);

	sysid_qsys_0 : component niosII_system_sysid_qsys_0
		port map (
			clock    => up_clocks_0_sys_clk_clk,                                              --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                             --         reset.reset_n
			readdata => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	timer_0 : component niosII_system_timer_0
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                   --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                                   --   irq.irq
		);

	jtag_uart_0 : component niosII_system_jtag_uart_0
		port map (
			clk            => up_clocks_0_sys_clk_clk,                                                      --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                     --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                                      --               irq.irq
		);

	sdram_0 : component niosII_system_sdram_0
		port map (
			clk            => up_clocks_0_sys_clk_clk,                                        --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                       -- reset.reset_n
			az_addr        => sdram_0_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_0_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_0_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_0_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_0_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => sdram_0_wire_addr,                                              --  wire.export
			zs_ba          => sdram_0_wire_ba,                                                --      .export
			zs_cas_n       => sdram_0_wire_cas_n,                                             --      .export
			zs_cke         => sdram_0_wire_cke,                                               --      .export
			zs_cs_n        => sdram_0_wire_cs_n,                                              --      .export
			zs_dq          => sdram_0_wire_dq,                                                --      .export
			zs_dqm         => sdram_0_wire_dqm,                                               --      .export
			zs_ras_n       => sdram_0_wire_ras_n,                                             --      .export
			zs_we_n        => sdram_0_wire_we_n                                               --      .export
		);

	sram_0 : component niosII_system_sram_0
		port map (
			clk           => up_clocks_0_sys_clk_clk,                                               --        clock_reset.clk
			reset         => rst_controller_reset_out_reset,                                        --  clock_reset_reset.reset
			SRAM_DQ       => sram_0_external_interface_DQ,                                          -- external_interface.export
			SRAM_ADDR     => sram_0_external_interface_ADDR,                                        --                   .export
			SRAM_LB_N     => sram_0_external_interface_LB_N,                                        --                   .export
			SRAM_UB_N     => sram_0_external_interface_UB_N,                                        --                   .export
			SRAM_CE_N     => sram_0_external_interface_CE_N,                                        --                   .export
			SRAM_OE_N     => sram_0_external_interface_OE_N,                                        --                   .export
			SRAM_WE_N     => sram_0_external_interface_WE_N,                                        --                   .export
			address       => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address,       --  avalon_sram_slave.address
			byteenable    => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,    --                   .byteenable
			read          => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read,          --                   .read
			write         => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write,         --                   .write
			writedata     => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,     --                   .writedata
			readdata      => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,      --                   .readdata
			readdatavalid => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid  --                   .readdatavalid
		);

	gate_timer : component niosII_system_gate_timer
		port map (
			clk        => up_clocks_0_sys_clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			address    => gate_timer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => gate_timer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => gate_timer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => gate_timer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => gate_timer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                                      --   irq.irq
		);

	audio_0 : component niosII_system_audio_0
		port map (
			clk                          => up_clocks_0_sys_clk_clk,            --                 clock_reset.clk
			reset                        => rst_controller_001_reset_out_reset, --           clock_reset_reset.reset
			from_adc_left_channel_ready  => open,                               --  avalon_left_channel_source.ready
			from_adc_left_channel_data   => open,                               --                            .data
			from_adc_left_channel_valid  => open,                               --                            .valid
			from_adc_right_channel_ready => open,                               -- avalon_right_channel_source.ready
			from_adc_right_channel_data  => open,                               --                            .data
			from_adc_right_channel_valid => open,                               --                            .valid
			to_dac_left_channel_data     => synthesizer_0_audio_data,           --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => synthesizer_0_audio_valid,          --                            .valid
			to_dac_left_channel_ready    => synthesizer_0_audio_ready,          --                            .ready
			to_dac_right_channel_data    => open,                               --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => open,                               --                            .valid
			to_dac_right_channel_ready   => open,                               --                            .ready
			AUD_ADCDAT                   => audio_0_external_interface_ADCDAT,  --          external_interface.export
			AUD_ADCLRCK                  => audio_0_external_interface_ADCLRCK, --                            .export
			AUD_BCLK                     => audio_0_external_interface_BCLK,    --                            .export
			AUD_DACDAT                   => audio_0_external_interface_DACDAT,  --                            .export
			AUD_DACLRCK                  => audio_0_external_interface_DACLRCK  --                            .export
		);

	audio_and_video_config_0 : component niosII_system_audio_and_video_config_0
		port map (
			clk         => up_clocks_0_sys_clk_clk,                                                                    --            clock_reset.clk
			reset       => nios2_qsys_0_jtag_debug_module_reset_reset,                                                 --      clock_reset_reset.reset
			address     => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address,     -- avalon_av_config_slave.address
			byteenable  => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable,  --                       .byteenable
			read        => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read,        --                       .read
			write       => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write,       --                       .write
			writedata   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata,   --                       .writedata
			readdata    => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata,    --                       .readdata
			waitrequest => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_and_video_config_0_external_interface_SDAT,                                           --     external_interface.export
			I2C_SCLK    => audio_and_video_config_0_external_interface_SCLK                                            --                       .export
		);

	up_clocks_0 : component niosII_system_up_clocks_0
		port map (
			CLOCK_50    => clk_clk,                            --       clk_in_primary.clk
			reset       => rst_controller_002_reset_out_reset, -- clk_in_primary_reset.reset
			sys_clk     => up_clocks_0_sys_clk_clk,            --              sys_clk.clk
			sys_reset_n => up_clocks_0_sys_clk_reset_reset_n,  --        sys_clk_reset.reset_n
			SDRAM_CLK   => up_clocks_0_sdram_clk_clk,          --            sdram_clk.clk
			CLOCK_27    => clk_1_clk_in_clk,                   --     clk_in_secondary.clk
			AUD_CLK     => up_clocks_0_audio_clk_clk           --            audio_clk.clk
		);

	synthesizer_0 : component niosII_system_synthesizer_0
		port map (
			reset_n                    => nios2_qsys_0_jtag_debug_module_reset_reset_ports_inv,                      --        reset.reset_n
			avs_writedata_voice_select => synthesizer_0_voice_select_translator_avalon_anti_slave_0_writedata,       -- voice_select.writedata
			avs_write_n_voice_select   => synthesizer_0_voice_select_translator_avalon_anti_slave_0_write_ports_inv, --             .write_n
			aso_ready_audio_in         => synthesizer_0_audio_ready,                                                 --        audio.ready
			aso_data_audio_out         => synthesizer_0_audio_data,                                                  --             .data
			aso_valid_audio_out        => synthesizer_0_audio_valid,                                                 --             .valid
			csi_clk50M                 => up_clocks_0_sys_clk_clk,                                                   -- clock_sink_1.clk
			csi_clk32k                 => up_clocks_0_sys_clk_clk                                                    -- clock_sink_2.clk
		);

	spi_0 : component niosII_system_spi_0
		port map (
			clk           => up_clocks_0_sys_clk_clk,                                               --              clk.clk
			reset_n       => nios2_qsys_0_jtag_debug_module_reset_reset_ports_inv,                  --            reset.reset_n
			data_from_cpu => spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata,       -- spi_control_port.writedata
			data_to_cpu   => spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata,        --                 .readdata
			mem_addr      => spi_0_spi_control_port_translator_avalon_anti_slave_0_address,         --                 .address
			read_n        => spi_0_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv,  --                 .read_n
			spi_select    => spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect,      --                 .chipselect
			write_n       => spi_0_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver3_irq,                                              --              irq.irq
			MISO          => spi_0_external_MISO,                                                   --         external.export
			MOSI          => spi_0_external_MOSI,                                                   --                 .export
			SCLK          => spi_0_external_SCLK,                                                   --                 .export
			SS_n          => spi_0_external_SS_n                                                    --                 .export
		);

	nios2_qsys_0_instruction_master_translator : component niosII_system_nios2_qsys_0_instruction_master_translator
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                            --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     --                     reset.reset
			uav_address       => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => nios2_qsys_0_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => nios2_qsys_0_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read           => nios2_qsys_0_instruction_master_read,                                               --                          .read
			av_readdata       => nios2_qsys_0_instruction_master_readdata                                            --                          .readdata
		);

	nios2_qsys_0_data_master_translator : component niosII_system_nios2_qsys_0_data_master_translator
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                     --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                              --                     reset.reset
			uav_address       => nios2_qsys_0_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => nios2_qsys_0_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => nios2_qsys_0_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable     => nios2_qsys_0_data_master_byteenable,                                         --                          .byteenable
			av_read           => nios2_qsys_0_data_master_read,                                               --                          .read
			av_readdata       => nios2_qsys_0_data_master_readdata,                                           --                          .readdata
			av_write          => nios2_qsys_0_data_master_write,                                              --                          .write
			av_writedata      => nios2_qsys_0_data_master_writedata,                                          --                          .writedata
			av_debugaccess    => nios2_qsys_0_data_master_debugaccess                                         --                          .debugaccess
		);

	nios2_qsys_0_jtag_debug_module_translator : component niosii_system_nios2_qsys_0_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                                   --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer      => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_byteenable         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_debugaccess        => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_read               => open,                                                                                      --              (terminated)
			av_beginbursttransfer => open,                                                                                      --              (terminated)
			av_burstcount         => open,                                                                                      --              (terminated)
			av_readdatavalid      => '0',                                                                                       --              (terminated)
			av_waitrequest        => '0',                                                                                       --              (terminated)
			av_writebyteenable    => open,                                                                                      --              (terminated)
			av_lock               => open,                                                                                      --              (terminated)
			av_clken              => open,                                                                                      --              (terminated)
			uav_clken             => '0',                                                                                       --              (terminated)
			av_outputenable       => open                                                                                       --              (terminated)
		);

	onchip_memory2_0_s1_translator : component niosii_system_onchip_memory2_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 12,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                        --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => onchip_memory2_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => onchip_memory2_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable         => onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect         => onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken              => onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read               => open,                                                                           --              (terminated)
			av_begintransfer      => open,                                                                           --              (terminated)
			av_beginbursttransfer => open,                                                                           --              (terminated)
			av_burstcount         => open,                                                                           --              (terminated)
			av_readdatavalid      => '0',                                                                            --              (terminated)
			av_waitrequest        => '0',                                                                            --              (terminated)
			av_writebyteenable    => open,                                                                           --              (terminated)
			av_lock               => open,                                                                           --              (terminated)
			uav_clken             => '0',                                                                            --              (terminated)
			av_debugaccess        => open,                                                                           --              (terminated)
			av_outputenable       => open                                                                            --              (terminated)
		);

	sdram_0_s1_translator : component niosii_system_sdram_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                               --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => sdram_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => sdram_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => sdram_0_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => sdram_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => sdram_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable         => sdram_0_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid      => sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest        => sdram_0_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect         => sdram_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer      => open,                                                                  --              (terminated)
			av_beginbursttransfer => open,                                                                  --              (terminated)
			av_burstcount         => open,                                                                  --              (terminated)
			av_writebyteenable    => open,                                                                  --              (terminated)
			av_lock               => open,                                                                  --              (terminated)
			av_clken              => open,                                                                  --              (terminated)
			uav_clken             => '0',                                                                   --              (terminated)
			av_debugaccess        => open,                                                                  --              (terminated)
			av_outputenable       => open                                                                   --              (terminated)
		);

	sram_0_avalon_sram_slave_translator : component niosii_system_sram_0_avalon_sram_slave_translator
		generic map (
			AV_ADDRESS_W                   => 18,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                             --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                      --                    reset.reset
			uav_address           => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable         => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid      => sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_begintransfer      => open,                                                                                --              (terminated)
			av_beginbursttransfer => open,                                                                                --              (terminated)
			av_burstcount         => open,                                                                                --              (terminated)
			av_waitrequest        => '0',                                                                                 --              (terminated)
			av_writebyteenable    => open,                                                                                --              (terminated)
			av_lock               => open,                                                                                --              (terminated)
			av_chipselect         => open,                                                                                --              (terminated)
			av_clken              => open,                                                                                --              (terminated)
			uav_clken             => '0',                                                                                 --              (terminated)
			av_debugaccess        => open,                                                                                --              (terminated)
			av_outputenable       => open                                                                                 --              (terminated)
		);

	audio_and_video_config_0_avalon_av_config_slave_translator : component niosii_system_audio_and_video_config_0_avalon_av_config_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                                                    --                      clk.clk
			reset                 => nios2_qsys_0_jtag_debug_module_reset_reset,                                                                 --                    reset.reset
			uav_address           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest        => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer      => open,                                                                                                       --              (terminated)
			av_beginbursttransfer => open,                                                                                                       --              (terminated)
			av_burstcount         => open,                                                                                                       --              (terminated)
			av_readdatavalid      => '0',                                                                                                        --              (terminated)
			av_writebyteenable    => open,                                                                                                       --              (terminated)
			av_lock               => open,                                                                                                       --              (terminated)
			av_chipselect         => open,                                                                                                       --              (terminated)
			av_clken              => open,                                                                                                       --              (terminated)
			uav_clken             => '0',                                                                                                        --              (terminated)
			av_debugaccess        => open,                                                                                                       --              (terminated)
			av_outputenable       => open                                                                                                        --              (terminated)
		);

	synthesizer_0_voice_select_translator : component niosii_system_synthesizer_0_voice_select_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                               --                      clk.clk
			reset                 => nios2_qsys_0_jtag_debug_module_reset_reset,                                            --                    reset.reset
			uav_address           => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_write              => synthesizer_0_voice_select_translator_avalon_anti_slave_0_write,                       --      avalon_anti_slave_0.write
			av_writedata          => synthesizer_0_voice_select_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_address            => open,                                                                                  --              (terminated)
			av_read               => open,                                                                                  --              (terminated)
			av_readdata           => "11011110101011011101111010101101",                                                    --              (terminated)
			av_begintransfer      => open,                                                                                  --              (terminated)
			av_beginbursttransfer => open,                                                                                  --              (terminated)
			av_burstcount         => open,                                                                                  --              (terminated)
			av_byteenable         => open,                                                                                  --              (terminated)
			av_readdatavalid      => '0',                                                                                   --              (terminated)
			av_waitrequest        => '0',                                                                                   --              (terminated)
			av_writebyteenable    => open,                                                                                  --              (terminated)
			av_lock               => open,                                                                                  --              (terminated)
			av_chipselect         => open,                                                                                  --              (terminated)
			av_clken              => open,                                                                                  --              (terminated)
			uav_clken             => '0',                                                                                   --              (terminated)
			av_debugaccess        => open,                                                                                  --              (terminated)
			av_outputenable       => open                                                                                   --              (terminated)
		);

	spi_0_spi_control_port_translator : component niosii_system_spi_0_spi_control_port_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                           --                      clk.clk
			reset                 => nios2_qsys_0_jtag_debug_module_reset_reset,                                        --                    reset.reset
			uav_address           => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => spi_0_spi_control_port_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => spi_0_spi_control_port_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => spi_0_spi_control_port_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer      => open,                                                                              --              (terminated)
			av_beginbursttransfer => open,                                                                              --              (terminated)
			av_burstcount         => open,                                                                              --              (terminated)
			av_byteenable         => open,                                                                              --              (terminated)
			av_readdatavalid      => '0',                                                                               --              (terminated)
			av_waitrequest        => '0',                                                                               --              (terminated)
			av_writebyteenable    => open,                                                                              --              (terminated)
			av_lock               => open,                                                                              --              (terminated)
			av_clken              => open,                                                                              --              (terminated)
			uav_clken             => '0',                                                                               --              (terminated)
			av_debugaccess        => open,                                                                              --              (terminated)
			av_outputenable       => open                                                                               --              (terminated)
		);

	sysid_qsys_0_control_slave_translator : component niosii_system_synthesizer_0_voice_select_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                               --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                        --                    reset.reset
			uav_address           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata           => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write              => open,                                                                                  --              (terminated)
			av_read               => open,                                                                                  --              (terminated)
			av_writedata          => open,                                                                                  --              (terminated)
			av_begintransfer      => open,                                                                                  --              (terminated)
			av_beginbursttransfer => open,                                                                                  --              (terminated)
			av_burstcount         => open,                                                                                  --              (terminated)
			av_byteenable         => open,                                                                                  --              (terminated)
			av_readdatavalid      => '0',                                                                                   --              (terminated)
			av_waitrequest        => '0',                                                                                   --              (terminated)
			av_writebyteenable    => open,                                                                                  --              (terminated)
			av_lock               => open,                                                                                  --              (terminated)
			av_chipselect         => open,                                                                                  --              (terminated)
			av_clken              => open,                                                                                  --              (terminated)
			uav_clken             => '0',                                                                                   --              (terminated)
			av_debugaccess        => open,                                                                                  --              (terminated)
			av_outputenable       => open                                                                                   --              (terminated)
		);

	timer_0_s1_translator : component niosii_system_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                               --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => timer_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read               => open,                                                                  --              (terminated)
			av_begintransfer      => open,                                                                  --              (terminated)
			av_beginbursttransfer => open,                                                                  --              (terminated)
			av_burstcount         => open,                                                                  --              (terminated)
			av_byteenable         => open,                                                                  --              (terminated)
			av_readdatavalid      => '0',                                                                   --              (terminated)
			av_waitrequest        => '0',                                                                   --              (terminated)
			av_writebyteenable    => open,                                                                  --              (terminated)
			av_lock               => open,                                                                  --              (terminated)
			av_clken              => open,                                                                  --              (terminated)
			uav_clken             => '0',                                                                   --              (terminated)
			av_debugaccess        => open,                                                                  --              (terminated)
			av_outputenable       => open                                                                   --              (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator : component niosii_system_jtag_uart_0_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                                  --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                                           --                    reset.reset
			uav_address           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read               => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata           => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest        => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect         => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer      => open,                                                                                     --              (terminated)
			av_beginbursttransfer => open,                                                                                     --              (terminated)
			av_burstcount         => open,                                                                                     --              (terminated)
			av_byteenable         => open,                                                                                     --              (terminated)
			av_readdatavalid      => '0',                                                                                      --              (terminated)
			av_writebyteenable    => open,                                                                                     --              (terminated)
			av_lock               => open,                                                                                     --              (terminated)
			av_clken              => open,                                                                                     --              (terminated)
			uav_clken             => '0',                                                                                      --              (terminated)
			av_debugaccess        => open,                                                                                     --              (terminated)
			av_outputenable       => open                                                                                      --              (terminated)
		);

	gate_timer_s1_translator : component niosii_system_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                                                  --                      clk.clk
			reset                 => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address           => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount        => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read              => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write             => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest       => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid     => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable        => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata          => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata         => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock              => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess       => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address            => gate_timer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write              => gate_timer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata           => gate_timer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata          => gate_timer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect         => gate_timer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read               => open,                                                                     --              (terminated)
			av_begintransfer      => open,                                                                     --              (terminated)
			av_beginbursttransfer => open,                                                                     --              (terminated)
			av_burstcount         => open,                                                                     --              (terminated)
			av_byteenable         => open,                                                                     --              (terminated)
			av_readdatavalid      => '0',                                                                      --              (terminated)
			av_waitrequest        => '0',                                                                      --              (terminated)
			av_writebyteenable    => open,                                                                     --              (terminated)
			av_lock               => open,                                                                     --              (terminated)
			av_clken              => open,                                                                     --              (terminated)
			uav_clken             => '0',                                                                      --              (terminated)
			av_debugaccess        => open,                                                                     --              (terminated)
			av_outputenable       => open                                                                      --              (terminated)
		);

	nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent : component niosII_system_nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => up_clocks_0_sys_clk_clk,                                                                     --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			av_address       => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => rsp_xbar_mux_src_valid,                                                                      --        rp.valid
			rp_data          => rsp_xbar_mux_src_data,                                                                       --          .data
			rp_channel       => rsp_xbar_mux_src_channel,                                                                    --          .channel
			rp_startofpacket => rsp_xbar_mux_src_startofpacket,                                                              --          .startofpacket
			rp_endofpacket   => rsp_xbar_mux_src_endofpacket,                                                                --          .endofpacket
			rp_ready         => rsp_xbar_mux_src_ready                                                                       --          .ready
		);

	nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent : component niosII_system_nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => up_clocks_0_sys_clk_clk,                                                              --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			av_address       => nios2_qsys_0_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => rsp_xbar_mux_001_src_valid,                                                           --        rp.valid
			rp_data          => rsp_xbar_mux_001_src_data,                                                            --          .data
			rp_channel       => rsp_xbar_mux_001_src_channel,                                                         --          .channel
			rp_startofpacket => rsp_xbar_mux_001_src_startofpacket,                                                   --          .startofpacket
			rp_endofpacket   => rsp_xbar_mux_001_src_endofpacket,                                                     --          .endofpacket
			rp_ready         => rsp_xbar_mux_001_src_ready                                                            --          .ready
		);

	nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                              --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                              --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                               --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                        --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                            --                .channel
			rf_sink_ready           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent : component niosII_system_onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                               --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                               --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                                --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                         --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                             --                .channel
			rf_sink_ready           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent : component niosII_system_sdram_0_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                     --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                     --                .valid
			cp_data                 => burst_adapter_source0_data,                                                      --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                               --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                   --                .channel
			rf_sink_ready           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent : component niosII_system_sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                --       clk_reset.reset
			m0_address              => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                               --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                               --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                                --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                         --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                             --                .channel
			rf_sink_ready           => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                -- clk_reset.reset
			in_data           => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent : component niosII_system_audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                                              --             clk.clk
			reset                   => nios2_qsys_0_jtag_debug_module_reset_reset,                                                                           --       clk_reset.reset
			m0_address              => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                                                           --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                                                           --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                                                            --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                                                     --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                                                         --                .channel
			rf_sink_ready           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                                              --       clk.clk
			reset             => nios2_qsys_0_jtag_debug_module_reset_reset,                                                                           -- clk_reset.reset
			in_data           => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent : component niosII_system_synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                         --             clk.clk
			reset                   => nios2_qsys_0_jtag_debug_module_reset_reset,                                                      --       clk_reset.reset
			m0_address              => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_005_src_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_005_src_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_mux_005_src_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_005_src_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_005_src_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_005_src_channel,                                                                    --                .channel
			rf_sink_ready           => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                         --       clk.clk
			reset             => nios2_qsys_0_jtag_debug_module_reset_reset,                                                      -- clk_reset.reset
			in_data           => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	spi_0_spi_control_port_translator_avalon_universal_slave_0_agent : component niosII_system_spi_0_spi_control_port_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                     --             clk.clk
			reset                   => nios2_qsys_0_jtag_debug_module_reset_reset,                                                  --       clk_reset.reset
			m0_address              => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_006_src_ready,                                                                  --              cp.ready
			cp_valid                => cmd_xbar_mux_006_src_valid,                                                                  --                .valid
			cp_data                 => cmd_xbar_mux_006_src_data,                                                                   --                .data
			cp_startofpacket        => cmd_xbar_mux_006_src_startofpacket,                                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_006_src_endofpacket,                                                            --                .endofpacket
			cp_channel              => cmd_xbar_mux_006_src_channel,                                                                --                .channel
			rf_sink_ready           => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                     --       clk.clk
			reset             => nios2_qsys_0_jtag_debug_module_reset_reset,                                                  -- clk_reset.reset
			in_data           => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent : component niosII_system_sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                  --       clk_reset.reset
			m0_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                                 --                .channel
			rf_sink_ready           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component niosII_system_timer_0_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                                 --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component niosII_system_jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                                                    --                .channel
			rf_sink_ready           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	gate_timer_s1_translator_avalon_universal_slave_0_agent : component niosII_system_gate_timer_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => up_clocks_0_sys_clk_clk,                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => gate_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src10_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src10_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_001_src10_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src10_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src10_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src10_channel,                                                   --                .channel
			rf_sink_ready           => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => gate_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosII_system_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => up_clocks_0_sys_clk_clk,                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => gate_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => gate_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	addr_router : component niosII_system_addr_router
		port map (
			sink_ready         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                       --       src.ready
			src_valid          => addr_router_src_valid,                                                                       --          .valid
			src_data           => addr_router_src_data,                                                                        --          .data
			src_channel        => addr_router_src_channel,                                                                     --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                  --          .endofpacket
		);

	addr_router_001 : component niosII_system_addr_router_001
		port map (
			sink_ready         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                            --       src.ready
			src_valid          => addr_router_001_src_valid,                                                            --          .valid
			src_data           => addr_router_001_src_data,                                                             --          .data
			src_channel        => addr_router_001_src_channel,                                                          --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                       --          .endofpacket
		);

	id_router : component niosII_system_id_router
		port map (
			sink_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                       --       src.ready
			src_valid          => id_router_src_valid,                                                                       --          .valid
			src_data           => id_router_src_data,                                                                        --          .data
			src_channel        => id_router_src_channel,                                                                     --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                  --          .endofpacket
		);

	id_router_001 : component niosII_system_id_router
		port map (
			sink_ready         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                        --       src.ready
			src_valid          => id_router_001_src_valid,                                                        --          .valid
			src_data           => id_router_001_src_data,                                                         --          .data
			src_channel        => id_router_001_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                   --          .endofpacket
		);

	id_router_002 : component niosII_system_id_router_002
		port map (
			sink_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                               --       src.ready
			src_valid          => id_router_002_src_valid,                                               --          .valid
			src_data           => id_router_002_src_data,                                                --          .data
			src_channel        => id_router_002_src_channel,                                             --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                          --          .endofpacket
		);

	id_router_003 : component niosII_system_id_router_002
		port map (
			sink_ready         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                             --       src.ready
			src_valid          => id_router_003_src_valid,                                                             --          .valid
			src_data           => id_router_003_src_data,                                                              --          .data
			src_channel        => id_router_003_src_channel,                                                           --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                        --          .endofpacket
		);

	id_router_004 : component niosII_system_id_router
		port map (
			sink_ready         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                                    --       clk.clk
			reset              => nios2_qsys_0_jtag_debug_module_reset_reset,                                                                 -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                                    --       src.ready
			src_valid          => id_router_004_src_valid,                                                                                    --          .valid
			src_data           => id_router_004_src_data,                                                                                     --          .data
			src_channel        => id_router_004_src_channel,                                                                                  --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                                            --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                                               --          .endofpacket
		);

	id_router_005 : component niosII_system_id_router
		port map (
			sink_ready         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => synthesizer_0_voice_select_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                               --       clk.clk
			reset              => nios2_qsys_0_jtag_debug_module_reset_reset,                                            -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                               --       src.ready
			src_valid          => id_router_005_src_valid,                                                               --          .valid
			src_data           => id_router_005_src_data,                                                                --          .data
			src_channel        => id_router_005_src_channel,                                                             --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                          --          .endofpacket
		);

	id_router_006 : component niosII_system_id_router
		port map (
			sink_ready         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                           --       clk.clk
			reset              => nios2_qsys_0_jtag_debug_module_reset_reset,                                        -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                           --       src.ready
			src_valid          => id_router_006_src_valid,                                                           --          .valid
			src_data           => id_router_006_src_data,                                                            --          .data
			src_channel        => id_router_006_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                      --          .endofpacket
		);

	id_router_007 : component niosII_system_id_router_007
		port map (
			sink_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                               --       src.ready
			src_valid          => id_router_007_src_valid,                                                               --          .valid
			src_data           => id_router_007_src_data,                                                                --          .data
			src_channel        => id_router_007_src_channel,                                                             --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                          --          .endofpacket
		);

	id_router_008 : component niosII_system_id_router_007
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                               --       src.ready
			src_valid          => id_router_008_src_valid,                                               --          .valid
			src_data           => id_router_008_src_data,                                                --          .data
			src_channel        => id_router_008_src_channel,                                             --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                          --          .endofpacket
		);

	id_router_009 : component niosII_system_id_router_007
		port map (
			sink_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                                  --       src.ready
			src_valid          => id_router_009_src_valid,                                                                  --          .valid
			src_data           => id_router_009_src_data,                                                                   --          .data
			src_channel        => id_router_009_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                             --          .endofpacket
		);

	id_router_010 : component niosII_system_id_router_007
		port map (
			sink_ready         => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => gate_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => up_clocks_0_sys_clk_clk,                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                  --       src.ready
			src_valid          => id_router_010_src_valid,                                                  --          .valid
			src_data           => id_router_010_src_data,                                                   --          .data
			src_channel        => id_router_010_src_channel,                                                --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                             --          .endofpacket
		);

	burst_adapter : component niosII_system_burst_adapter
		port map (
			clk                   => up_clocks_0_sys_clk_clk,             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component niosII_system_burst_adapter
		port map (
			clk                   => up_clocks_0_sys_clk_clk,                 --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => width_adapter_002_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_002_src_data,              --          .data
			sink0_channel         => width_adapter_002_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_002_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_002_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_002_src_ready,             --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	rst_controller : component niosII_system_rst_controller
		port map (
			reset_in0 => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1 => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk       => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset_out => rst_controller_reset_out_reset              -- reset_out.reset
		);

	rst_controller_001 : component niosII_system_rst_controller_001
		port map (
			reset_in0 => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk       => up_clocks_0_sys_clk_clk,            --       clk.clk
			reset_out => rst_controller_001_reset_out_reset  -- reset_out.reset
		);

	rst_controller_002 : component niosII_system_rst_controller_001
		port map (
			reset_in0 => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in0.reset
			clk       => clk_clk,                                    --       clk.clk
			reset_out => rst_controller_002_reset_out_reset          -- reset_out.reset
		);

	cmd_xbar_demux : component niosII_system_cmd_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_src4_endofpacket,   --          .endofpacket
			src5_ready         => cmd_xbar_demux_src5_ready,         --      src5.ready
			src5_valid         => cmd_xbar_demux_src5_valid,         --          .valid
			src5_data          => cmd_xbar_demux_src5_data,          --          .data
			src5_channel       => cmd_xbar_demux_src5_channel,       --          .channel
			src5_startofpacket => cmd_xbar_demux_src5_startofpacket, --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_src5_endofpacket,   --          .endofpacket
			src6_ready         => cmd_xbar_demux_src6_ready,         --      src6.ready
			src6_valid         => cmd_xbar_demux_src6_valid,         --          .valid
			src6_data          => cmd_xbar_demux_src6_data,          --          .data
			src6_channel       => cmd_xbar_demux_src6_channel,       --          .channel
			src6_startofpacket => cmd_xbar_demux_src6_startofpacket, --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_src6_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component niosII_system_cmd_xbar_demux_001
		port map (
			clk                 => up_clocks_0_sys_clk_clk,                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			sink_ready          => addr_router_001_src_ready,              --      sink.ready
			sink_channel        => addr_router_001_src_channel,            --          .channel
			sink_data           => addr_router_001_src_data,               --          .data
			sink_startofpacket  => addr_router_001_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_001_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_001_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset               => nios2_qsys_0_jtag_debug_module_reset_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,                 --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,                 --          .valid
			src_data            => cmd_xbar_mux_004_src_data,                  --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,               --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,         --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,           --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src4_ready,                  --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src4_valid,                  --          .valid
			sink0_channel       => cmd_xbar_demux_src4_channel,                --          .channel
			sink0_data          => cmd_xbar_demux_src4_data,                   --          .data
			sink0_startofpacket => cmd_xbar_demux_src4_startofpacket,          --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src4_endofpacket,            --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src4_ready,              --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src4_valid,              --          .valid
			sink1_channel       => cmd_xbar_demux_001_src4_channel,            --          .channel
			sink1_data          => cmd_xbar_demux_001_src4_data,               --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src4_startofpacket,      --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src4_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_005 : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset               => nios2_qsys_0_jtag_debug_module_reset_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_005_src_ready,                 --       src.ready
			src_valid           => cmd_xbar_mux_005_src_valid,                 --          .valid
			src_data            => cmd_xbar_mux_005_src_data,                  --          .data
			src_channel         => cmd_xbar_mux_005_src_channel,               --          .channel
			src_startofpacket   => cmd_xbar_mux_005_src_startofpacket,         --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_005_src_endofpacket,           --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src5_ready,                  --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src5_valid,                  --          .valid
			sink0_channel       => cmd_xbar_demux_src5_channel,                --          .channel
			sink0_data          => cmd_xbar_demux_src5_data,                   --          .data
			sink0_startofpacket => cmd_xbar_demux_src5_startofpacket,          --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src5_endofpacket,            --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src5_ready,              --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src5_valid,              --          .valid
			sink1_channel       => cmd_xbar_demux_001_src5_channel,            --          .channel
			sink1_data          => cmd_xbar_demux_001_src5_data,               --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src5_startofpacket,      --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src5_endofpacket         --          .endofpacket
		);

	cmd_xbar_mux_006 : component niosII_system_cmd_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset               => nios2_qsys_0_jtag_debug_module_reset_reset, -- clk_reset.reset
			src_ready           => cmd_xbar_mux_006_src_ready,                 --       src.ready
			src_valid           => cmd_xbar_mux_006_src_valid,                 --          .valid
			src_data            => cmd_xbar_mux_006_src_data,                  --          .data
			src_channel         => cmd_xbar_mux_006_src_channel,               --          .channel
			src_startofpacket   => cmd_xbar_mux_006_src_startofpacket,         --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_006_src_endofpacket,           --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src6_ready,                  --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src6_valid,                  --          .valid
			sink0_channel       => cmd_xbar_demux_src6_channel,                --          .channel
			sink0_data          => cmd_xbar_demux_src6_data,                   --          .data
			sink0_startofpacket => cmd_xbar_demux_src6_startofpacket,          --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src6_endofpacket,            --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src6_ready,              --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src6_valid,              --          .valid
			sink1_channel       => cmd_xbar_demux_001_src6_channel,            --          .channel
			sink1_data          => cmd_xbar_demux_001_src6_data,               --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src6_startofpacket,      --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src6_endofpacket         --          .endofpacket
		);

	rsp_xbar_demux : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_003_src_ready,           --      sink.ready
			sink_channel       => width_adapter_003_src_channel,         --          .channel
			sink_data          => width_adapter_003_src_data,            --          .data
			sink_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_003_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset              => nios2_qsys_0_jtag_debug_module_reset_reset, -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,                    --      sink.ready
			sink_channel       => id_router_004_src_channel,                  --          .channel
			sink_data          => id_router_004_src_data,                     --          .data
			sink_startofpacket => id_router_004_src_startofpacket,            --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,              --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,                    --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,              --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,              --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,               --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,            --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket,      --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,        --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,              --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,              --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,               --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,            --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket,      --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket         --          .endofpacket
		);

	rsp_xbar_demux_005 : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset              => nios2_qsys_0_jtag_debug_module_reset_reset, -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,                    --      sink.ready
			sink_channel       => id_router_005_src_channel,                  --          .channel
			sink_data          => id_router_005_src_data,                     --          .data
			sink_startofpacket => id_router_005_src_startofpacket,            --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,              --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,                    --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,              --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,              --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,               --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,            --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket,      --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,        --          .endofpacket
			src1_ready         => rsp_xbar_demux_005_src1_ready,              --      src1.ready
			src1_valid         => rsp_xbar_demux_005_src1_valid,              --          .valid
			src1_data          => rsp_xbar_demux_005_src1_data,               --          .data
			src1_channel       => rsp_xbar_demux_005_src1_channel,            --          .channel
			src1_startofpacket => rsp_xbar_demux_005_src1_startofpacket,      --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_005_src1_endofpacket         --          .endofpacket
		);

	rsp_xbar_demux_006 : component niosII_system_rsp_xbar_demux
		port map (
			clk                => up_clocks_0_sys_clk_clk,                    --       clk.clk
			reset              => nios2_qsys_0_jtag_debug_module_reset_reset, -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,                    --      sink.ready
			sink_channel       => id_router_006_src_channel,                  --          .channel
			sink_data          => id_router_006_src_data,                     --          .data
			sink_startofpacket => id_router_006_src_startofpacket,            --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,              --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,                    --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,              --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,              --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,               --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,            --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket,      --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,        --          .endofpacket
			src1_ready         => rsp_xbar_demux_006_src1_ready,              --      src1.ready
			src1_valid         => rsp_xbar_demux_006_src1_valid,              --          .valid
			src1_data          => rsp_xbar_demux_006_src1_data,               --          .data
			src1_channel       => rsp_xbar_demux_006_src1_channel,            --          .channel
			src1_startofpacket => rsp_xbar_demux_006_src1_startofpacket,      --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_006_src1_endofpacket         --          .endofpacket
		);

	rsp_xbar_demux_007 : component niosII_system_rsp_xbar_demux_007
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component niosII_system_rsp_xbar_demux_007
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component niosII_system_rsp_xbar_demux_007
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component niosII_system_rsp_xbar_demux_007
		port map (
			clk                => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component niosII_system_rsp_xbar_mux
		port map (
			clk                 => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component niosII_system_rsp_xbar_mux_001
		port map (
			clk                  => up_clocks_0_sys_clk_clk,               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src1_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src1_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src1_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src1_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src1_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src1_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src1_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src1_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src1_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src1_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src1_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src1_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src1_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src1_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src1_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src1_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component niosII_system_width_adapter
		port map (
			clk               => up_clocks_0_sys_clk_clk,            --       clk.clk
			reset             => rst_controller_reset_out_reset,     -- clk_reset.reset
			in_valid          => cmd_xbar_mux_002_src_valid,         --      sink.valid
			in_channel        => cmd_xbar_mux_002_src_channel,       --          .channel
			in_startofpacket  => cmd_xbar_mux_002_src_startofpacket, --          .startofpacket
			in_endofpacket    => cmd_xbar_mux_002_src_endofpacket,   --          .endofpacket
			in_ready          => cmd_xbar_mux_002_src_ready,         --          .ready
			in_data           => cmd_xbar_mux_002_src_data,          --          .data
			out_endofpacket   => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data          => width_adapter_src_data,             --          .data
			out_channel       => width_adapter_src_channel,          --          .channel
			out_valid         => width_adapter_src_valid,            --          .valid
			out_ready         => width_adapter_src_ready,            --          .ready
			out_startofpacket => width_adapter_src_startofpacket     --          .startofpacket
		);

	width_adapter_001 : component niosII_system_width_adapter_001
		port map (
			clk               => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset             => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid          => id_router_002_src_valid,             --      sink.valid
			in_channel        => id_router_002_src_channel,           --          .channel
			in_startofpacket  => id_router_002_src_startofpacket,     --          .startofpacket
			in_endofpacket    => id_router_002_src_endofpacket,       --          .endofpacket
			in_ready          => id_router_002_src_ready,             --          .ready
			in_data           => id_router_002_src_data,              --          .data
			out_endofpacket   => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data          => width_adapter_001_src_data,          --          .data
			out_channel       => width_adapter_001_src_channel,       --          .channel
			out_valid         => width_adapter_001_src_valid,         --          .valid
			out_ready         => width_adapter_001_src_ready,         --          .ready
			out_startofpacket => width_adapter_001_src_startofpacket  --          .startofpacket
		);

	width_adapter_002 : component niosII_system_width_adapter
		port map (
			clk               => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset             => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid          => cmd_xbar_mux_003_src_valid,          --      sink.valid
			in_channel        => cmd_xbar_mux_003_src_channel,        --          .channel
			in_startofpacket  => cmd_xbar_mux_003_src_startofpacket,  --          .startofpacket
			in_endofpacket    => cmd_xbar_mux_003_src_endofpacket,    --          .endofpacket
			in_ready          => cmd_xbar_mux_003_src_ready,          --          .ready
			in_data           => cmd_xbar_mux_003_src_data,           --          .data
			out_endofpacket   => width_adapter_002_src_endofpacket,   --       src.endofpacket
			out_data          => width_adapter_002_src_data,          --          .data
			out_channel       => width_adapter_002_src_channel,       --          .channel
			out_valid         => width_adapter_002_src_valid,         --          .valid
			out_ready         => width_adapter_002_src_ready,         --          .ready
			out_startofpacket => width_adapter_002_src_startofpacket  --          .startofpacket
		);

	width_adapter_003 : component niosII_system_width_adapter_001
		port map (
			clk               => up_clocks_0_sys_clk_clk,             --       clk.clk
			reset             => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid          => id_router_003_src_valid,             --      sink.valid
			in_channel        => id_router_003_src_channel,           --          .channel
			in_startofpacket  => id_router_003_src_startofpacket,     --          .startofpacket
			in_endofpacket    => id_router_003_src_endofpacket,       --          .endofpacket
			in_ready          => id_router_003_src_ready,             --          .ready
			in_data           => id_router_003_src_data,              --          .data
			out_endofpacket   => width_adapter_003_src_endofpacket,   --       src.endofpacket
			out_data          => width_adapter_003_src_data,          --          .data
			out_channel       => width_adapter_003_src_channel,       --          .channel
			out_valid         => width_adapter_003_src_valid,         --          .valid
			out_ready         => width_adapter_003_src_ready,         --          .ready
			out_startofpacket => width_adapter_003_src_startofpacket  --          .startofpacket
		);

	irq_mapper : component niosII_system_irq_mapper
		port map (
			clk           => up_clocks_0_sys_clk_clk,        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_qsys_0_d_irq_irq          --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	nios2_qsys_0_jtag_debug_module_reset_reset_ports_inv <= not nios2_qsys_0_jtag_debug_module_reset_reset;

	sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_write;

	sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_read;

	sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_byteenable;

	synthesizer_0_voice_select_translator_avalon_anti_slave_0_write_ports_inv <= not synthesizer_0_voice_select_translator_avalon_anti_slave_0_write;

	spi_0_spi_control_port_translator_avalon_anti_slave_0_write_ports_inv <= not spi_0_spi_control_port_translator_avalon_anti_slave_0_write;

	spi_0_spi_control_port_translator_avalon_anti_slave_0_read_ports_inv <= not spi_0_spi_control_port_translator_avalon_anti_slave_0_read;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	gate_timer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not gate_timer_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of niosII_system
