// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.1sp1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H $/0WM_53O0)^OT0T(HRF=BY=_M"XP0731VL[Y'[_\,B1^"NO+5"%   
HP>G.(D-H<;3/FE 8PT90<O@VR;]Z?&9],MZ+(A>-TN.*WLNL'C%)?0  
HS]GD+R8MF;)L203-]C"]SFM[L3F?[3;4<O 5/O,*V,+RRBT$J'COE   
HX#%$/O)_%+T6>?0ZQW/_O--I%SQ^WM*ZT$!L,M_@)[J  :-ULI%X9   
H^="E!3-)5CJA#+EEF.CJF7JFO*AH:^]?7V[WS?<EI2 DVG',L-WIT   
`pragma protect encoding=(enctype="uuencode",bytes=12608       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@_%FK<GYD23SYZLCSJ:/^CBN0\O+*6EE%@<\P:H+<F<X 
@:#ILH\!.-U3^>;LT?R94U9*(C.UWG3Z" *6I'A3;HRX 
@!B6HV7V 0!ES#P )-*Y90+LO]CT[^ L WE GF'4P@8H 
@:$T ;P^<8+_('P'/JL^S&?D+/(CI+(G543V GM3 T9  
@N[LTD3S6O)U]7]<%X-BB]]>P068AED\ 7TXN8.UUB)0 
@T57SJN6LB%(\YK\@0W29T*8/E *D#>-C0?X$T. ZK;P 
@&O_4F$8,'P7S*LG\@'BUEO-ONYI/.L/!*0.L*U.Q9=( 
@YV74P\9W#ONR[M>*$)75K6D7Z76#R_GZ!>B&+FT4.Q@ 
@^%H7QM[Z4IAIMEDISZKY.F(K]^&HU6HB8.=^XXW4JQ( 
@NZ&OAI@@1<HG$!\G@R_5+*3%->$&!)"!28G&,<"UI0\ 
@]UL/!@8JKS#-@@C\T1?1?X,?#]JT1IV4KQ"@4F0WBQ4 
@0+CF"BX_6(.NRHF,#0D3N;/3PRUF)-?9JJ^2J*1(,M( 
@=7,C?V"GGO/8;5BUY9ZB^IZ=ZJ8_67F"7/S_G$\RJD0 
@Y#DU%EH77@4EZ#]V/NZSHMNYF.CQ&(34L,@LIDV7=0( 
@PN0"\;ZL<19! )5M->Y.8$ .+WG<;*9LAZ]644?01W8 
@PC+TB4*2YJ^&&O26YEC"J52_S^>-P"*DRRUR"CG -\T 
@P^RT]@S\EW:WY.5B\QE(+6F+NK"3<=^9EV\U/0626-  
@8XKV'W0:0.K+OQ]QB@>B\5T,H04XO,-3%Z+^+V$*AJ\ 
@!K;$4*9AX ]@:]K!)(UOAN6ZBV49G[NZBM(X:A\U@+$ 
@:-R#;^/'&.LX_7 K^\8VFNS66O ?<-T!UI1<E*:'!%( 
@^ A[8L0%PC JB=/F[J_YR"9SL:DO#SQJ1XB:4_Z1VVD 
@EDR5U+3;PKHY82";LDWND 4D3V6!%Z5@1-'-8 ( Y4\ 
@J@(?Q2W#ZAL?F@P@FFX;H*M_[A'4;,=B7T6^&]: C'0 
@E!>U_+F/;AD.'U"#[ G<<?'U_]';Y9>D]-4L-QM3: @ 
@G:?,GF(RWZE32CN&>WOC1AH'*1E5H_=.%&8=YY!VQ[4 
@R#E,>G.&#G!"K75<(U&<,K13DT[;UI OZ4<#!!J!U!, 
@MDHJ5O[V@J*F^&;HE\?(RKTD2 [O*9OQ@PLU7 AI5R8 
@C&/5=EE?ACAH*!4P<S^+PW'2LPM$\N++I.Y2DEB [-D 
@"$3%ZO>(MTSQYO&DK7H]Q7#P.B.U#'N6R>S[W'P ,U8 
@[":^#?9@-QZ3F%02Q 7&8/W!!0M?>/5%?QVIF>UI908 
@AJ%*X3T9V_E%GRL'2Q!O!/E7E(FL:BQ'<T7O]%5J+UH 
@)Y@R5#0BH_TTC!5%95 I56#ROF WX%]*:,I;]+49%PH 
@0FQC!.DC$",H&ES@&<7=V[X9N7Y+BQOEMS1C@FSV)@\ 
@7Z6%GJIQQ(L^U8!'!M6\&1>GSM*Y,[(P^51,39NL?_8 
@;?\55:F7Z_#J!FCCW=K/%_!><P:WY _KH:I?D,Q#V>0 
@]$-!,'%][')NQ)"\*,A.>10TFL53#N=7I[04+;.7[J@ 
@_)@?.">8YP,T.\V)6#*BC=N!:;>*Z)NT,4K+#NF6H'H 
@SW%@MGQ:L%<M!1T6Y:+@"/AVD_K]Q*UT?733!39FYY0 
@4\US_L]Q<7(ZD=0E_8G0?:A:XG<^P&[J-P%L[[JX5>L 
@2(J?YZ&R-$\W-46(H>7]ZP'A:#;2'P.>M,HR&3@VEBT 
@Q&H.]>.M2XI//4;K1FUZT H;J[$[JK4!X7#9<6!E5F, 
@5*F$)S)YZR_$.U4=H[#:U>XN%LD^\)J=!3U:5[0?F:$ 
@-<!V__*@B&5M,O1"[/%TX"\M*:%C1;P0Z% 8E3#>5+\ 
@P,0WA9!!:A([E$A'/J:MN2FU,@?Q)1 YO?(\QE2C)Q, 
@@2F_C;OZ5><_**P9?1-AQ*%BY8"KZTI;T&_TVS:Z%J8 
@LXH/BK+OF5<A#].^>3B5EBXYUE]-DUO\I(D&\E+T95T 
@4-9D(7\0^0_M5/]U>?$F:BGC6#E-0F>B9)HAX'-VO'< 
@VP4<.S9U0.ZM_P6R^_\H'](-"CH;?1>,1W696[$?X+D 
@0@QFT2E)[]M5@_4,BI==4?)MJOAFZ\ J;K)![FQ02YP 
@:G"<CT_1U2RFO>00Y#0<12Z,($BZ'1*;,365PEAY3@, 
@#&$8\Z&2J 14VVLPG 1Q;FR&%K;\0S<O%=6$=5;! 1D 
@:-&9#NCBI@4T).0_O-:U)'BN=0(#  @@8 !_A:BV?J0 
@;9W@V)\;PF5<*)XL_B);X[K(>G^\YJ)AWQ:;VL7N5FX 
@>(O1N&7_GH5),7 DDI;RPN;O90EWJZ@K 7!DVURI1*$ 
@L287Y[V'=:':*11!_TXF&%4_&!!4JP]2[RY_T^K7L   
@= #TXA\P"=YIOEJ6T4;7QR8S1'U$W/535%(<YB!OL3$ 
@41*^?X)FA^0"L)FCJ=G#5F^<6Y/Q/K+1OV06U4U2AX@ 
@!H8A(.<_T>M+GOKBZMP]W'S!4"S.R%>1 ,>P6.1>[G$ 
@<XGGB X[P;8FO@LN'3HC*()4L.YU5K 9C@[K4&;3>GL 
@.\@I#)AYY9-*N$%>9!]CR"BTW(Z%@WMJ4P0X)_7T"N\ 
@!+8K'3Y&9>;*%>+2JI9P)H&L$!1+BVS!QT+:?\0;L:P 
@E9,/:#MJY%_F-//,0L@X/%J5#HNNQ8WH=J*2=*;X%_T 
@HJ^D V1TR;VK(_A#:JOG"1LR4&8U0 $D)3V"M\53@4D 
@QIY>ZM(-$&V5?3Y01UINJ6Z&,'$C"%+;.@,M?E5++HT 
@8$=VM[8Y81K\6LW"F;PO%F8<9:(Z47%J/:7?G#T9RR4 
@_W<H;UE#OX4UJRR:W&_Q?69TEF-J<@TAEF[?.\I] TT 
@+6,Z+(.9&): M-"4TB'#Z)A@T)?G-^JT0G UEF<GP.$ 
@)Q^JOI35T'"K*EN(* ^WYB]@8R:QC;X<2+!3\-J6*G@ 
@S/HRHO'DX5>7VKU(,%Z9C[7,)O (._8O\@H3_XPS.*$ 
@F\LZ&6)-\J.6MIB1]K3X.@0IINCRXKC6;!B*8SCZ5:4 
@W5KF,MZMQQXGK&RC*G*\N[OW/5N9RWU.);=E8. 3DE( 
@X\&WM@@ED]25W+YX7(F:N19&CD3J%'O]9[DATB1';DL 
@7/S2*( QJP[_&_:JM>? '";-:(/L[DH,7$U.+WM*29D 
@(,V:FA-DAK#F_$J_7IRK;ICT\ G5$3,3&V)F_G>NQQ4 
@+1V^CART$:[:-OEB^0^AN!A< &.U"&*-2)$TV5_9J?$ 
@S\*+)2.,:DM#1[?U*M-VM,A\P5V''[2Q8;\9;>(ZMEX 
@@H820:RB0)G,A*GZ)REK!D_3HT3W"?M!3KX%6(AKU]8 
@>UT>> E?Y0V-$4PMCUCO.#-K[..0(+QSA'4]#1B(?;@ 
@V--F@8BRRN_[?O=L*[UX7K"%2"#HJ$9B?U'-.$&DA+8 
@M)9IP@+N/N/B/7DQQKI7=7; _G->5JA4 =&2$11@E&< 
@EYO#E'WAWUK\F*59WY2'A:-Z3&+O) -$I*Z;8GNDGW$ 
@IQ'F$&:JT]#%I*_)XI10E7E!+H24-W(-0:PR6 H@4DP 
@.!8;#U"X .AFL&XQX!/7S%@BJID2Z(6 LB-481+02IX 
@#S-Q<'%LGY77?CJB \D,L135AG[?@\>\>./Z#G-G,/L 
@R&)6,YKN4^]SD'Q:EP_K<=:)<5CK!T$0*UO3^O*\L*0 
@1,5\+5Z&^M3+9VSJS-$$J2</&:*V%B[#\@L[5\RY@RT 
@_1=)WTBG6'95I,B@5_K0Y L UTKM1Y]JNQG\DTOA<$4 
@LR[V-0KAHRM3=F1YZK31,N&$4 #_SM7Y_61G)._+\"T 
@90X'Z5G=XH%)"T.;[-!I:%C7CSF!4MAHW-#5@G O#=D 
@=1-8'!2?PZH%=5004797KI==4&9T*D^0/GDR_<-"I.L 
@7U:JVH&$6^47Q7__<C\H)IG&#5KGP\THWS*04 IYS3D 
@)U(F=D,#71LZ>LV<('8^!E+-3FQN0E6(OCPUG:&>X%\ 
@$+I"4)Z^H#DZ:6\OOH"!2R!^UU6>@!PI+/KP&9FV!*D 
@[UVXL2-3I&1RQ^O$.;+MGU%%05J[R/P\2E$%X\1I4P@ 
@"^'-42)M#%E5>7N6EJ,N6()4LD[,@&:_#7+X\=-@V2H 
@WP%O,^VF6)\Z;#:,N//C,A193M7V"&'&3D:%\B$9-X8 
@^H%57*7I 9W=EEZ=)FOAU+N!CJ5;2%3DV,.'&>ISYYP 
@U\W%T-\I%I>%URTY?;$>W@J^+GS$7DQE*$DA4]O$P&4 
@;Q"+AFKPTB3O#G$K+)_SHYTIA[U?R*!.WG0/CYY5R5@ 
@ 0UMXZ"^K":DL^3*E"![-I/>1X*JT@Y34J-1TH U<?  
@>R<]MEEL2U"0DJO]>T':_$%@IY]YT7PRV!,\<L(D\RX 
@Q!OVH+*+,0D1/@TF2VU99.X7X<N.$^@)3S D#][)S^, 
@V&?2U1E!AO<?^XZEN=-A$]%!=)MQ8O1 "YJH9GT_M0L 
@D1TR*#GV3NW8> %YZ@43ZK'%V:(0 DG)@]=3O.=*?Z$ 
@NZOEQ-SWZ3>25RA0!7C\]% ?SK/CC'$20=];2+['DI0 
@CUEP?93$F"9*$(];AJY&*QWD,#9I1ROW1X_6M% )8DL 
@'""SZ-GT+ S\=P8(WR:EX<Y!5-23OW.1$ZH+I*KZAFL 
@F7R4O$G(S:729M;.-PFQ9C?0&U7U%3*66R$1@63W3S, 
@(AE&G#FV-OL"FUT%Q^Z+$<[?W:ZZDVG&;4#/ -\\SS\ 
@0[^MZZ!R@+DX=:0 JI/HIQ^#/;2OA:E\)NFW!UJX.94 
@8?8/8T+?CE Y($QL2P(P?N1J%2?L5>)B(^[S ZUO[_L 
@F_"2 DO)=LY2&^&0+ R'$9G4+8K+QBM(3DF *2QC/:4 
@6ABHS ?7?RAM+]]B#@M,MT0B)5P[6Q\G#M78:IT$&CH 
@@(S&!FGX>%W_8*=0KO0PY-CT2/VFWX'0>F8NN_-V$]@ 
@T=E,$&]G^.]>N&<.XD8\W%=^FBX.U0B33O_U\U8%,?@ 
@HD^?_PN2R^UZ$A$H-M#/L+:1[.^R.DK?"CCM:W;D]Y4 
@![$"#F!HB^%5$BS:<A[U5R-),!^'0DHL,HOV,[)2NB8 
@E$GF8$Y\M+O7F6.$CJ&1N&A_S+S[.AN8[/K+B=;.D?\ 
@N8N M!:OK#YZZ8(]KU'/4K+4>)6:[)XI;FF7>MB9^"0 
@!RF:APUKA' 'F3'1/Q"9^QHRIA+E8=Z7L,Z,9DT5VIL 
@'R[P) ZB,FO;T%$TYU7KVG:;1?US"E;,'L5LQ-T'%[8 
@MDTU[4",3YY-;RZ[&L^EX^T4J"F)HN3R55E::VQP43$ 
@U!"!HN'"2X2(U6K&;RV]7"QQHTQ;Q_,H%3,QWJ[..)( 
@GAIFPH*V"26WB2QJXZGX-D=Y=/KX#OPO= SUBG<Q-R, 
@LO+JIV8?K/3=Q %FD;HGVZ'+!+0"8!%"HA,_*Y4+&>\ 
@T= )$NUZ()7E)J?,BJ@6G2Z\U%-AK?DQA[4/@.7J#U  
@:73M.46#![P#;B3Z)_5$6K%*"HR/6N["['Y)=5/[DQP 
@)GO7#P@@6J7-3.%:VX'1/3-W"P$[V_T"BCZ=)PR3@Q, 
@!W=:X)PLF7%,,87O?3.[H1J!9D,Z3GW+."Q=\<@Z2A, 
@UF!W?E<SXA+?@=2S7S%Y.\=9Z/Q+E>IK'Z^#6ERA,Q0 
@NF [ZKU( 2-)Z08<N<LY6N ;97N2R/2]@^$6%S<DJ@, 
@[0!B[QI?])II@A.@3J;6/$*;#]H7W@QM@EF8K&F>\/L 
@F)68+\/;1SC*\OJTB$3B RESJ!D>F@XL->N_%G\R7QX 
@+.+"86M^BH=M^*5D4:)9@KD=4Q ).JHVR0#>ZP?'[0@ 
@C_B8B5F7EMI':+N>JS1V/A>FV2%&4,34>0685W:TTTL 
@/]^'?)6HGZH!I:&-XAURXKKK&UT-3:]9-C@2&HTMS*\ 
@KB1PL6[Y#<D4;^$Y;VI6-M8=Z@:"IS<8HG!]5Y2G_WT 
@F11GPW0L36'K:EH2Z7+IEHWV4B+DQ-&XI[GWSVSK@ P 
@ +7&=?49NZOR%S[ '5$WZ$L_8O#_9WNF43=$]Y\)>B$ 
@<LHB,T\<&D;@7?]RI_;-,*IW 1#M#38.7&,X' )M.:H 
@.(EU'M,FL8+J/<71D8^VB.<!X ?'BGM=0 <!><>RX]$ 
@NOK)A"<\O^-H#3NMKXM3E:)_[=+*\RV-E&,<D=S1TQ< 
@TXPG-C3F\I0VJ4;9\ ^/TU$DDL/).C<5IX6.A].*PPP 
@W3H0G,3SL9'&35Z!'7:FUV-#^4G[C>XS8@#S96LTS9< 
@7@OH=6-)JZ3NY2/L&%T;9PO4[Z?C0>U;+"?(%%X%52L 
@$6Z(*T8[#<,('WC^W;\V": 0+V09D&<L%HK*\9)W:UT 
@9%)KYI]&A125RE5.WMPL6FGA?*N)EP\ EC3/('O,0)< 
@U<0)Z1M#1UC(G=U;"FE/WR6ES\Y3(!<D+*,(N HHFIL 
@AD;NF%5)R0-M4.DVEL&[@0VK">_(AA90_9Z*514+YV\ 
@SG^DJ%N/<AX1;/I2CHD#^S6Y<QYP><'W+)PFEUF4".D 
@B2CB[L]&1&#1=#=!H2@[N)?+2RX9>C#H-H3Z19[L(SD 
@)TS^QL2U+8?[T^ 0HW'N4-]W-K'WN4F,H&Z;+5;O#*\ 
@92SL41""L1F@N"%4UX(-OJ\8=[X->*+4I'7>-CQ;)), 
@+!_2()?+9U%+_2?244[ B3\G?O0G6V0E#G(_ED7P)<8 
@JUD7SYK 0$:[@PKCP)6"M E%!<GS;#U+]Y*1Q90%U:L 
@3@P:Z-<TE',Q: 9B/F</RIK J;T3]44)?V1P797)9@\ 
@V#.\<+)Z1^'%\<A.'?A*PH+NK!Z]7@6Z A754RN8R*T 
@O-N#.IS)3@)8ULN1!O=\T4EZD[;3S^-LGUVHGA%_?+P 
@;S.Y,UOV+*2GR31A?,OQY #(BSGX1'!LE $ S2UC*ZP 
@#6M;$)B6@SXY&(Y7@XF<%<1/M1 )-:)IAV>1DDVW6F8 
@1B7S]PFG6Y>'2M:A7N4^3.M"PWA'># Y!WZEH%^+0TH 
@ U1P56!&QG,)="%WWRNI;E9<ZVW$I#VD$<#;6J:^ZC< 
@C66C/1B.^+7G)=P/#FU4]>53<H0!L!\+\\\;Z!/[7ET 
@$=C4P.LM%S!@PP2,C$T#"A'"216^)#5E#PU ""R]B(8 
@!#!-S+EX.6[T5VS"&Y#)9?5;A'ZC$!I(C9GALP*D3XT 
@BMS+@2=&M)'RHU7#9J-KV6L?)UL5Y4@N)R[0LO!: $@ 
@MQ96L+U!,OK0B@E'!_WD<K,,=;MGB<.[WN_,[K"N/ X 
@N@==,NF'01K:",\&-O8'SI?09EJ4"]NGQZXQ=+;-6^4 
@CLNK!6\:<_S5G &Q!!DD?<[;U!2,@"('[-G*WU(3!-@ 
@UI1M?S?U\,&\C6P&Q>!1@CZA$1QV(!^,[\>LF;/57DX 
@+WG7K2.ZA'U76E\V6%)GI2;DA8(.^F)20VTLTS4."]$ 
@>O;'?1MU$GC(@T2Q5J'*_:)-XTAZB/'\!I9XEA@(:?L 
@9N%.;[8Q^Q\L+D])C?Y)SZHJA?[-FAD6!%,OU1L$]Q< 
@Q72(V3D# 9\'_148H[/>@=SP0,7+-*&=AEB\[%!JFY0 
@%K/>/2T8& >!B:+VIH>*&^D%D\8-):&1$X@70++)KEL 
@%Y"EFE&"^N[X1@5AM?)D4\A=Q]XX.3;LB:Q??IF(\%4 
@,@Y/=JH0N+F'TW)K .2)=\>#@'D**Z[)\8!R[?KL 3@ 
@-1D.L*V4DC#O[K-02+!G=\^E)X;7:S.K*M0)*D=JXY$ 
@I1EAHC5:'>PG^L@U-TR.M3HT*&8<"AZ[D;ZPO.YQWB8 
@T"!R.R<T54PBT/F VHGH@D<!R]-2 ZCJ9*9++,?2N@0 
@@I:B ##/LXXV99K8FK&SG>+%Z!.KJ(@H'GDV-E6^_@  
@[@$6U"C0&F.>-\>]0#A9LUJAQ4UJN0V?=,[KX'W WU( 
@N!AD&T^P#7%)L^6$B_*X5RF<R>*'VQD@'>,13\ZHS $ 
@CT2%@<#+48!_DJIE"JXK9)1[@B:QBNV(2_EQG6GO@T4 
@2W.D4 K<NINI@9R"863C3!T)H9@W>.K080ZX.2A(<\L 
@O2ND;D3V/W-]_5%?^K#:PS4R@F>"K$P8^<#<)9/2I#P 
@>+CXNV  W"EM-]IE@S@\R W(LL@MD3,J=F.\>I(00(@ 
@=FE0B$H!*>GA?*,%B^!G]GF3>[>4_O)B]C&_+&1\GYH 
@ X*AS+SURKJG:XF,[GV=0N^:,Y$\I6/,3?.2>Z"%&EX 
@P.=U1A9"NY/DP=491JO0VB:7Z_B\.&!B(?+G-WFCV6L 
@[=ZE@D3HU-H5##I>.@DXRVZ9WT*UC,1TP2]][9/?/D0 
@D[8<6-!E?963Q[!; KW9[J];N>K&;'+ZKE0)@RJ4U#( 
@;,A>NH?D\M[R<$V]@CW<Q'P]9O442,:L787"?/9]3-$ 
@4K-HA6OW_J-4QCHK+V752&R]AZ F(TIY:77:DLRA>AD 
@8F+D]'A$N<(\>W9C ?:2] :[KM2]?5[:2\@NC:OH2/$ 
@W?*=LEE;D%VYM@Y[KTD\8W*L6[3M+5S!--@,^\:NX), 
@C"M3>SDL!$+.:F?(K2 [)1V-LP-WU5MU;5_T:>W-A+4 
@VOLI6(I+]4U\T]%%2;WKF./Q2;G'F9+_QQ]-I.T4QA0 
@-"*\24N)TY ?X1WEJ?^S%M2B%VKS+6V?\H2)"T&*#<H 
@4?5#K3=-?C7[DX$9P JCR);T>A_@NI,V J3.SI8U 5< 
@UW;AI0?3(/*%9!?H1H&1?WC>%# DXU@.NKZ#W'SQDN< 
@DI :LPX7!18E"@BS,D'3' 8(%]!G]138;5O5F-IH)<< 
@H6S+W>XN;,IM<D />FU5C!807554$8.2Y;4I?^_4_7< 
@X_W\"8*><R3)08;06U;%5WOG!;OQJP#5II3X6,<*AWH 
@2*S[>A)!4)68BAILC7)+;1_"GX]2\M+E+H!8=?<'N,L 
@)_@(//FQ&\X"\IBN(*"Y^"X3R! B)>%M9WTP?&2A)$( 
@8*01+]00^Z*GBZ..H8EPH^[V%8I0\GUV_!7A2P<Q_WP 
@,,JQ,<8>1VA&L-JY2UD5+:_5T1+A51HV'KV@W>/Y5I0 
@BE>G-ID0A$T:=7V/8]IJMVY88X$@RSP!!M5:D9LN+,@ 
@?[/TT]JC@IJ944>GQ^\?0F':W8+^4F99N)?MB&-NW\$ 
@JS,3THPER54\>H<N->*X<&=\( WV.6BZ=R60LLP#T!H 
@$7Q^M?S,4A ,%=(;#Q8K#=S !HM2"!.!#L":GAOX["L 
@!CAU?088PBRP&?N X)Z^+LWQ$*N5'D!@+^ :D ;C(GX 
@[W1BI;N0J>%S?&AMO1(82WG2>V,C.66N9[A+6LT,TMP 
@& >F6V O3V=MZI !=#VCW_7-;]7>?"8.^S7R\+6.7PL 
@ H*H#[7>C/__6"I2'8/)_D[SZ6\'G#_,.>(G]&7R!^4 
@:?Q.4.7@X"@)_1%;XD@U(LHJ!-4+(/4OA;4?+W_"N 8 
@4$Q7U^6OQ+]]1FA?-CF,,Z)2%9[FOX--2E49&!8>.6, 
@%XG'Q7N"KUY3 =F?,O)WVPF8U(:(*=0(<*$. L)9HMT 
@?8J3^DJQ0;&JI298ME<.VD# _;!1K[MJPC-CK"D'+I4 
@QF<IC0MHUNRG/*&;B#\ZL1J+G0;0UFI]W5TR$7PM/&T 
@0C8SNI1]1=)TZ"L&Z6.XEZ?<1;@]7>CP8'EP*FE;8ML 
@@7SH1\UKZ7K=/BCW!GC0#&3&3T8Y\;>HU N)=7(_&O  
@6B'K]0C&!RP'<T"?#19!U"]92T@2#]V SAT1Q+U[<$8 
@#][CU^)Y)0C;H?2:\Y[AIXIU"![Q11L:CPZO0#MKT?0 
@R1MYN'FJ1G2(QHN[WLN1_PA CM3MK8\/"CH&C0A0'4\ 
@)_*,:P5L=N1<5X$N]-S_O-@_H%P%9&RUGJ#',GTZ$A0 
@=ED]OK8L2X$\XB0%O#N4Z'Y?72L-NWY<\JT,6& ZB@< 
@@\6L<"$T4I?K7Z@ W;>]Q<^<6-R_<!PVL)R/%3 =B1( 
@I;821 Z402B/E7!5]2BFXP19'\G=QCM73:*M,1*!22P 
@H7$#A7-F<J5%H_0:GK(/_<U3DKN3(YIC88/!&4I):T0 
@TE !/<7\;#(](V8=\KRS@N0.8MD@@]ZI&=$@A)V9S)( 
@XD!/[*DFU:3P-ZN_[/@L.=P&A1I:;&228+R$SC%)29H 
@-!)Y"J-#;3-KUSCXHHY[)XMRENXV;/ 8S].8] .EH1T 
@Y;59,20]%?'T@RA6)*CPUQJHPO=.5!/MQST4,8X_( , 
@[P?&8=SL]P,ZB<8ZO!&T[LP4C@IZ4)RRC?!%:N+A'<X 
@(OY3(M07%C"'FT-:8(N]?/!K5X&O ))Z+EO\K7^>RO@ 
@*UHW=199EKV,3M7+2(C57YFQ JOF^=I_% LV>VD<9(0 
@X/X1LXIL+5MF>9HP<Y#;\Z3OY9#(VCB*3#W.W8I&9[, 
@RF9JV88[M#0N9C8WI"0B9.M/B FGWBO^BN66!8L$9$< 
@UB:B9&)LL'.$)GS[[GWOD4Y<>S7:H0WW@'[?@BX/_L  
@%]U[M$@5,&DM\1^^05!5S4;@\7#0%R"-F)L(E*"Y&G< 
@-R^":!9JC%W_EH$RY66U6&HF93(1-!+9L%__7[=1J8  
@R_@_BYC\\5(UV_W <I80U\*,$,6_LKGN#\G3-JN\JM  
@#M%GMKO_/.AB[[Y=38E4V'R[=7>EPI$XI:O:N%@$-W  
@]X].-CU#^XI8\.-"R(PPKYNJ>9 4UV>\0:T=.H&*X), 
@*C(UM^Q)&6W\%^?M;<LGAGP\[AB.OV)5^ /1[U/Q:;0 
@?\@Z]!2'[$\*N)T=Y-#T?H0#'B1>D/8%OO[OR,FZQO8 
@6O0+SJC_O</EO03#*NO[ 87T+71&F<MP-8VM9)J$RI8 
@KW(P\^RTN'/N_>:U Q; BL"$)&9K&\!!,5;/J;4O-+$ 
@YL63_M8*EH.0%Z^-0KDH3&<78Z7-NOT!<&U@:3<,JNL 
@0;-=/QO2UEVZ?.)DG44-]L4EH!ISF^4Q?=K#5GD!Q\\ 
@^X%>V#!;J(O:,]&BUX):XV^QS6,2JG%1N4?:'S$94R@ 
@J9>98P<T<"+)L>I/KG/S9H^VE=%#_EY!"O@V$%L,(14 
@46!GV3R!;DBG</7/^URO+F,@W7^)ZTC1>,>'(U)@/QH 
@WE35 E(@*S4B%5>2:T.8%9<!E8M]BHP9"?(DA 4 IPD 
@4T/Z%C T A-.8_34XY OYZ%%VU3E7J^U?,2=1.F/1C8 
@J0Q#MFNITDHE5E[+AC]P]WR\'7P%Y.^FD!A=#H5-Z=0 
@Q1F<MB:'UKTK^FWZ>XCX%W]U^< !6K DS0^7=NRUQ=T 
@F,<<LB2!R#U"E,_N^@3:W;*\"K]+80@)$")Z#YRT()T 
@+Y%M@FQ)[<,]L+VID;THI'0UXA+(;IYQ2HFV'[U3#&( 
@]KS],56M#',^1O2* X<]-:71ZLV#UM/HU1(!3H%,?\  
@\>"2%M,6!_]H2UE\"\0"-"E:WS=LVA*%59//=#C+HXX 
@@M44-1MKOMU$#9V@(J^$U,67M\X.9S]'46^[U6XEU]X 
@@JGO_)%Z>I@M(C'@H9/HCT8[%HM)&L(A%FISOY;Q4TL 
@5BO=1\4FPHT9+5!29UW11(@/U9E+QUA@O1=P/^U9V4T 
@KQ?3*(Z-<9^\,<^L U/1@72QV9:9['0QD]0EKI>%@B  
@/U)-[<SQ4F/VF3OB?27=%@X"LQHF-+B]=OE_9N#E]38 
@'?;]H+I/O)U+\VAYM'&'LX#)M#PT=P==CDP2@V>AM5\ 
@>D5E7L1Z1,?I*#5N2*J=46/#RSS*RAA>K-)VQG.IQ&@ 
@$&OH^\0;(EZ\O3-P6?GV](_02^]P[IEO<\:T/:%\L[  
@3M\;] 0AYKH+ +49BB16)G9A\H<(KCEOT=!L&K1B*2D 
@VM#A\C>IR>8ERJ4ZP'$?]VE9J5//X'$6AA(I=J.(#FT 
@75SQ^H-=H$84PN4B%C?;R7P# <\&S%</7!5J78<TZ80 
@"^ZFR'D%;I?%(*&0"]XLD9L/1K(?N=#+G[>GP@[*&20 
@)&%PE,KC\_DMA/%2CI-F\/(7ZL0AJIR;5$0U^ZY)@Z8 
@/N2[ VN:DC?^@ KFG)9J_T AW^0QL![//%KA.7R+Z:T 
@4@QGDSN6 @VWQVLZZ; K^U05 '\2Y!'YWC\"N3#047  
@ZBT)CC&_E/4#5[+M7I$B8F4LI5.>XL&5Y_= S0LQO\4 
@LC$FV[-E9DB\D#G8[.;K%N><56Y1RM1P!.A3[]4D"-D 
@G$<,#:Z?A=GT_5!+/I;QMR7!V1AWUG 4YNF0]S74X2H 
@( 34#5Z(6)97;NC/TM \2^M/\I>\>\^D.7)K;%-?X^L 
@*01ZJEW+;5-,LHC66KH([9H(S22WRSR)259V4Z_< KH 
@?@Y C\G@LN<<S$WBJM<I02:-1M"RVFE#$IC,$@0T>(D 
@R?RQ'*.S 3MBA>"SKG!IXK5/L'- Q$W0J6..SD65<@T 
@]&\5.155"=*7EP!\R"D,5;A[PD3\-F4_MHZK?'\QVU< 
@=3Y):G>JW6U$K$DF<H$TB/K.-2^';! KWL(V,3W73#L 
@YT-U(+?R3(+!Q']EJ)@MWI+9(_%F#/?./;#X3:QE@)$ 
@^;)MLH'JV$U?X*TNN#?M$P6B%>IO3M4"3N9VWE+D$54 
@6.P)P!D5YR+:D+5$R<!+ SZ;&F@4"W(H4]W>9GMK&=< 
@SEM.!%[X?*C?Y3\; #0Y00*NGEL^XQB D( V4T%I]]H 
@2ISNJN,H<32>6\O&Y:L%O[ -I>;K[_N55YU4@UD/Y&  
@V"A3RRC2V-Y%R5T#,SN;0,-+G&6:9",*'NIS6[C<N:L 
@-"=7GA\Y.K2]4C6]4BK9="\XYDJ5)ZH1E65;KO-+H$L 
@EON5-/H61S>!.KO3#X$PD&?].RB\*<U#Y"4C PT&Z<L 
@:EM@X4J+/'P8V'^<J]QNSD]:70 T=%-?6?<W.$785($ 
@(9^&4ZK/4KS -L6HIM2'!"U]1[BS0P@0V\N=K A6_PT 
@R*S)Q,AM+',MXE0S)",1>N\\;X%?M&YI)U:=FO!N./< 
@*02R8>X X5FRJ5D[ @,)(%-(#:-P4+MVO]8V'C74E@0 
@LEFF/I700LD6W7'L<_V?3?[;07_NKUZ9VR)5][C%-<, 
@X!",\K>R+I^QY/JM_&_WR191VE@(W8[QS4I"Q(9CPGD 
@5N$6! , 1&UJ;M4-NZIJQ=\B*:ETNA\<K!K &W$ZS]X 
@7C?[(])-!<):U^(D9[-KH2__QA14Q6(@8!OOV3X!2-T 
@\)M#BR?[ECP(Z?^M1/+$_<9'B_07HI \;Q\E'?^1Y"$ 
@]:6W@O%L$=:*Z2S[Z& Z7;VQP_)\#C4G4,W\]:-IM$< 
@E62I,\Y%X<0D 8.%Q[9H\2U\+;_O?4TIK"9C,YM][ 8 
@7OIOY"%P9[%VCF< _Y'_)E"3 \'SVAV\72W7/U?EM&H 
@PN%?;%\+:PR<2(HP7X2/4;/3 X/::@GN7M>N>$(LR,4 
@-E[O&JF&>NZKKL@/=#>,;-E*KXQ0Y(#;)U@#G*0HY]D 
@1_Y*Q=*Q5FSLS)Y3IH:@:JTR2XJ9@3P(*&E>&*+$D+L 
@D&G?@,?U[/12'6^)OHA;W!#*IXQ,8C^&JMQ6V'!H5L( 
@C.=KRT\ZHDQ)QN0? 8;E@@V>L=JKD7FXQNZ^QJ;?OB\ 
@&UFW2E B3[Q^DQ*JE^"#S%H 4.^5FMCQNC_7_UC;]CP 
@7H'OP-.:H%T.<^[XT7]33?*']AQC,WTE[0OL[S XF+P 
@WY6SEA8KH!;YWRNJIK4<G9%2T_WHU;P1TJ^JRH]B/%X 
@7/\@9SATH0Z,P>M=14.(E&*5:G.KK9 9J=(8Z(>%]:T 
@TSRE\<D?H(<846WZK)"<F3XG"HO6R#_Z;AW6Q:@AHMH 
@T5E"NUFY;M@1BK*%LR'ZH"W@$R0CEQ'D>,'#)FU!DM\ 
@\;P6'^R6E3Q3N<^,>ZK5/P9TM>- %'2/<PDC8A3H7QD 
@DZ"@<3"4HBGH &'8[$XH/"?%CTJ)0&^A6ASZJ35WQGL 
@7:!:>@1UMR[$$1N[*5JW+"NZEG/C'+/*)T@0Q^?XMS  
@$>NNJ4@OLP#\3")'P1A.X.)US7%GV1O".P',T)_S@[H 
@^#6\/B:$'$EMS"2$08XV7L/1.JIE$_2*Y8ZA&WA&M]< 
@-8#%&=E$'2UXHM]5-J9<W788JPXX9,,31B,=N^\YR#8 
@!;_VQIOLI!0S#J*@6ZJ^!0%<Y,Z+:VY@,'WA H(DZHX 
@YJ"P1EI<)O^O5PC3X@WA=,Q'O]H5B,!YZUR+R3MN$6X 
@'# /J%1+9&UEN\[$;8"Y1"4@C:6&+4'&=^^G9C=\1<4 
@&QG1ZT9Y\:4#Z%QH<G/@CFE@F,:":P5-%1&TDYK0.5  
@NH5,?&T9GQGUXGR"P[?T+& #1HOO<;Z*"0'2/@:E/Y< 
@;Q>B");Y/2#?\$$N<S-U*>>7QJW)2%-*@N "MSZX],\ 
@V+DBNL)*N:S#S\M6N"N_@&_SLHU9<;^G31@I=P;!SL8 
@-,2*:5K!B8\\ZAI@G.)AIQ_+\56E\CL0]2=L;J'$\<H 
@4EI#K]*;-MCI2%D0[#I;*UQX2,3N2'SI5'$(@P]5;,D 
@%Z+FMAD+?/'K'30$9@V9&M*K[7BRFQF8"Y5:4? #5E8 
@B"]2*CD3=2D0\@_+Q(%1K70_XW6]**FDX8Q.01![(#4 
@5.;%0$4*^8D0,K9HA4G/@I$FSU(?7L>7HB>WVN$7NJL 
@\:I=)J!15!/?M7C9##BX]=>THUUDN4Z)-N<-Q9[ )&D 
@NK#BD.B:-::!VAN[^G%?9X9WKY@+VENZ#PD?Q%H^XL4 
@.\\XR]K^R,]5 X*"2HMQ22$[NM3W8Z8\&X_XSV@+SJ( 
@"I,4T8G*_<;DHBW2*[)Q35Q+M@8'TTUE29N75OHI4R, 
@@V_]<0"_/57BOY!_XIO(./E$VA7I-E:]-W>%2V"@BEX 
@DKP< =?%B*4Z"D!+LSC+V;GEG7D:M-61'M3'E''DCO0 
@%L_LIL&M/VYVC,OFQ)@1\1>U;R0/U-\T(@)9C(-K"M@ 
@&T4 410MGK2=X'J+'L63'NNNIC]IL#!4634'"Z,Z2)@ 
@;A7V1^XW]6#5$H@J 1P1-"4RG<^%FJ,FY89]*K!4M<@ 
@T(>O+ 9$LVWS4A&EE^.MM#XK;&S+OJ?\BQV%\3!5=MP 
@)Y,8,=(3R/]Y]PJL^PQY2E=/#+A"HSJGJ:.^V)WV1B8 
@05FG":<,\Y%H$@I+("=5OL^GZ;ZK]_8'Z)+8AN7L&VT 
@\DF2&4.8QD<F5"9<AJQKWI(%SR7QB:(F!N/''A654GD 
@92;:%1S\0E-"7=_&=^S[UGK/=5?',MA2$DT'NI9X(6P 
@<P;75EC^G_HT$/V/W"3CRC5_4D3L;_5DWW\ )*DB=30 
@![C4&A7/:*FCQ,R_P>T!0A6@@GPO,!HK=C91%E5]DM8 
@S2]W@ZQB> '\9Y'3N0\;Z"H#)6I1];!;+RN<V\K7J%0 
@94Q(]I$7A[0I0+RL6-#Q.G*D.Z/U@+DKF)RR*,H+@0P 
@0;A^ASEZLG_;07I2;H%DTUY/>#AOE(SY\HI29+)[/-8 
@G1W'_C?"OGJFB;F$5@VCE(A-IHFD0;]A.)O%R U4E&  
@!I&QI@.JWGIMV7-!)SA8+W XUQV_KK4R#J&S+<WJ3O  
@DZI29=!^.J@_()&&8()V1[J-FVDM( BN1Y8ESO G%?, 
@\KB$0R8TUFZPXRU3,KYVQ73DP5;U'CE]U2<A_[/F8M@ 
@2#=<7?HJ(_*!C^+]22[GK#K=A:U*>NSN"+2DVT&NP@( 
@K(6VO( >$5?$XHXXN,B/TTA>-][C:&B%34OZ*,H2IMH 
@"; -4'[<:SU4#9( "VKPQ13WL$D1IAS >A4B&-,V/:\ 
@&<83GS_]RQ?OIN#LFAH]]K5J V';Y-@3#-_6KCA_MWP 
@- 7VZ"O])<C_C#1)PW6R"6EF^F=.ED6EH9@"H4G)>8P 
@A_N<JP/8)AGRKT0QL)<X/@(_J,X(T=TI 35QZ@$@XY$ 
@6-JT!:S>H;N*H $N7[/+@73%LW*G@YV>/BPBEL@L]ET 
@JJ$BJ^GW%)(!Q^!ET4N.J,CZG3Y^4Z4#]20N %G[2?( 
@9QAU*N[[@%=$5<U .YO@^('7O<<YG1]* (G2!T; =%@ 
@)T?VX8@8F<S\.7MH)=@%5%F (X>H]_@NK*P5\%?\,)< 
@A3)8E$TBTOBB<E8FGO:(Y2=[/:FAP;CB^1'XMN02XU8 
@A$@GH^W:7*TUMFDY2NKH)1H>Y>;,7$W0E!@N&+EE;8P 
@/CG"Y651E>%M"976FRI1VU2P32B=" WR(VT1.K**!MT 
@>O-=L>,\\GK<DCJX#!A049%"3 GI$T^W'=ZE+R0C%;8 
@8>Z.J()GQ!/=?8G&FNBK&P9%?.;+JDW=Z,N%IZ)CUG$ 
@QVO -/%.-ET19M)TYQ#[8ZQY/<C.E3>L6BP'_ ]6.>0 
@WO %E:-6_LXP<L$V2I';,MT&.=-G/CC;RCM-CI,-]/T 
@(W&AYVCDR!BB!EAECE"Q.,]IY8-PU9Z8 TC8G,+-H5< 
@]LUBI<_NU)QS*O/E2Q.#XQ[\"*F$#MXZ83Y=A 4D^_( 
@K<87^E_:L1@;WWQ/_A\24S:E(ZSO5Q(E;4J6=7 ]YO( 
@T'LPK;\.)+893^9,0>K<.(Y)>#Y]AA@M@^A7;'?MJ+  
@=V+&0@_0QKE\=MF$%.QV4@^1K6:E\J)6IXJBQ9GCYAH 
@V,>S.N$]=[-+;ZIF&EK#!=%)PGON>PTB$3)C)G+<D=D 
@V*X-T6D'><!6RY,?P29(\1=AYDP1V.=3E9]B>)E_&N$ 
@/5[#;XUV+[32#B _NY$\E/-Q?Y_.VQ S,K"NZ2%:IR( 
@_@(*DQ)D<N$/] A4ZJ._+XMFS2*-1B=$-:AW5@-V/3  
@$ ,"FM]4Q,%-B5"9)<6CF-+6T+^"!1FNM/D/M;G*_&@ 
@O^HQ-K+V2\0T=_YC[T08K-J8WWUW5I:]&"=E1^^I"(8 
@4LVJ.S04V:?^SOKW4XNJZ@3<*O"]+-(D<:3H=JU;P04 
@5Y^SLB%>:#"_7M$Y&A3I'4,N?@"I%3I$AC\;>TD]49, 
@=9$M<2$CH[1AR/&280,6VR[.N1\5BP/S'?;P6+)5E>H 
@B"SY%.G2/D,T"MXWS]=/XX7P2:;KZS-$ KV/1DF[2S\ 
@<+'$JF H/B_G!_T#IO8!?RSG3@ZB1T=J_&:=*LS_*B< 
@, ^!JW>^/$J6(U;*:ZC&VTG(H9OT\P9O+2>A79 "#UD 
03P\6@R(YP;QO<##>&?JO>0  
0,\&XS0U.I4X5J K#3-)ND0  
`pragma protect end_protected
