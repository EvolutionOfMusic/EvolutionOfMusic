library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package SynthesizerPackage is
    type PHASE_INCS is array(0 to 0) of std_logic_vector (31 downto 0);
    type LUT_ADDRESSES is array(0 to 0) of std_logic_vector (11 downto 0);	
    type WAVE_ARRAY is array(0 to 0) of std_logic_vector (15 downto 0);
    type MUX_INPUTS is array(95 downto 0) of LUT_ADDRESSES;
end package SynthesizerPackage;
