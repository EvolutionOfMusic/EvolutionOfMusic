// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.1sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
PQtMRF62fEjHgYtMIM/k+l/Qohi6oKQrDeq3tFmgKphKDc1ueehJJS3dAxoEvnvachDURwRzT+pX
k4cUgBaYxWe/eXPnDWxoQmU/B1c+BbVB86+qOKWWfgORsUJJLwDOqBYUz0/WF8SlD3+XTRNXfpbq
1G9C0QBSIuyyf2RravvslguT3KUtnTHmScq9ydahR3gPIPJOrMfsTHV2WySmOdx8l+vqVE9mVr5A
217VHBwSViB8cZP4QGcTa1laolc3k6h4lFEU1xWGZ5FGMe4go5blu8ZNkNzsDRuL1Ja5HlIJQ8z+
AwspbuDNIP9djCJR0UMY6O8mmiyzHBkywtOSOg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
4tv3sEhhWNdQ8U+cP1pQmfzF+Yhd7SqX9v+AsXsYdqglgX8W0sI4sYBXUlJg+W0hK5U/ONrc/1B4
ukridg+mBCW0qRegGxsKHspnITfmlqJOe0Qc4Xv1MGu3jDQKG1qbwiKjm+efD24T2eOzgi4Topiv
mHoSyiUSGuAThueSn0Ct83EW43hlgGABMU7kCeyDOK6rPQUQ7ljVm1UDhhepDHYzgyhVLtQHSDEa
ODKwRqKLWrtqORYE/jcenfVWGb+ZQT1Kn73FRZyjaRIvrCtkoyIcOudVX/9QYUDBO7kVTg/ngXvc
ANQ5ts3n99FeNyXBCV557tYuOdv4+Ay9lsnoWsAedqhvHffCu6Mshtr9S3JBjtnpLVOnZFBJDdYY
KZ5JTlB6SF7WkI5lw1Cr1ZhcAPSytaM6jifIOKxrtNlFk/Q8j8CWB3Nmy57GIbjn+/59GiVI8/d7
TJAcTBKdmIAAt0S5OT+oqMICM99NTUvTh7XFXL/wzIp+NpEi19N41WR3hvKuwdox/3DB9cTi+A3q
oEr96couFnTBXVCsmw01WSHj98ScyrH22vB3cDCwSlCFbkC1YYKlc1laijq1NH0dQvnFp8G2b7TL
tAhywLNzSad9LuSq7qMEe7Kl+GLIdOKAOi1KbBlspB0Wh8mOp9E/i8t06P89L28bR40Zxg5dLZ3E
1fC/kFeSy7hFg6/U6EO02wdJKqXxdmx8NZy/hs34tmfLXEurQdZjgV6VdOI0a4gnPs+qcGHHrm+e
Eca+sSFAT0oO/GYodESwdAc36b2uZIkOhDiUuh8dbVxBTcKmIhJgN9V5hu3M0jvXW2Al/vKMEi1S
/qDoVcY0OTUp78x2iKK/wWpQxQa0/NMLMafzYI69kYhgoUGZvdLB5V6a5KfFqAy18EXd7bSlW/8v
/oOTB4Ixrx1PtuYCHj2BKwr7iVyc1w9Hm88haG73qtvlyqQyG5BNEwUDVEMbMd0b5y2H1EmtJ4qv
4TkF74Lh7wTm5X4WxRHa+Bv5cFJNStOit7b1alz2gCD/N1JT6jkrtWWBfBHD7ulMIiwpybgXBkKn
OpNhl8/VX9jR2xXbSrjBDL3zW09y3lDuZmLKsmoJ2kQpDvNVt2EBM5dD/xTQk1XOfAjG3uzcof+y
HbDX5vpIFDgteyIggF84h2HI9mgmxwCYJmT93ZrHSiqaKNGoAyavMPdyHJGRz6imnNQybgaAzmcX
UWMZGdnkDvUlevz9XaPlrSo9Atod79TogV16t4kuOB/a2RkCQfxsIq7n1vH0ylRwE5Xm87hwj79S
LQBH/A8Ef1Ll8n/K9K2gX8rCB6mgDbgQj+4TJRJ53jslgVqnp98Ln0jLranfAL8LJp8Ay6qoArK+
qlUfeeZeil2pcTXntGCOy/eQcL23D897s5av3kIuTZD7zQMaLqXt3SBRVzdUIqg1CD3Xh+/2qcOg
zk9MfhDVquE42ZdduybY+MGFe8O7xOm4vyAV3jzmR92K3G9UbGbNP0nIe1yCWMt6tsu0814nedam
jRMliyDO9TQ4zzvBsWyzJpH1JxGXbef4rkyaPaMa0WIHG+Cd7AlETGNeClPa874ySL0BZHdrfchd
pOZgsGEa8XSfwsJdZ8536dRvtCazNWUPFFT/PA4ZPoSXUr/Nvh6HmDugWdbnriF6EmgOhlTm3Jy0
8CtO2YXIOGJKlI4EhXaQxQhv8YfE/QjOYj5Dr0IpZ6e/kpCrsZdDeuMp+ollEvFf0sXZ4ol/l03e
RIyIJ6voF8ZdT+CbAo6viWC9TGE1veneo1yRpVqm49I61qPL3bjHQ0lf3M4fLqQasssdwP1xrIWf
vGrZTX+XE/60RE4w0xsITw59IzH2zERGigIE/3hGpQBJCq8/CuSijCS3UeFo+MAqI1048wuQZIxq
lyeCLqvN9MWLy3I25eLXy2WE2fgpQoZX2W2jb734nf5ysiLVGjg6tOGl8uZSp+LGgfEbMUYVGfQr
Gz0txUHpFExpaMFLIsJrWOEwWqV2KI93P9/yjG2fNub/C2elXT1eBQtClcGIQpulbS+oknJPdAXk
34cALe412q6iAQ0kEQJDZHxVUduFVjrGcAS3g5Gq5B/y69Fkg+q8TnvrTQUHj7rvYWq3z5mJ7Otw
o/U4pHZVkT4t7oIhK2/ryTUV5P3gCKlBNIAGNUw9HAH8juCYjxVFwv/NU8mm/un//bWtD3akP7fG
1apTYcw1i55uMkMwHkN1TNV3VDqJ0r1qT3ag13bkmfxXq3k45bQ+YIWzdX7DDEr7G0tXrkr8/9DG
mqBovMvt1tRhqjJi9Q+udt2s5HBqijfy0yDfqDTm+vRulLerES/7PSkOMGVrljvBJbNsAz66iwYM
b1Si5xQCMuhCxa//ocY+d7IH9jI27gkiw9EsJcVGLblTa/Rgs99CKpqm26a5Os5uej6pptuhEWa3
Zi25NquMSCLbLS2AJNljxfXdBNFWfZDSfTQ9Lp2VF3wGjFQ1JP13JdBtiR4Hg3ZXIz+e7rvuikmp
PRMwZ3k9QSN7UmZjiV7s2RrZyV6ykGdho7NTgVPcRVT0epK3sqzo4PviSLXD0dRvX9ISKVdsYzv2
271OT9d9u1LwshswNFcqikXUN8xxeHVcvNkmQI22ew92Ccmt+RlyLIX2tZtkBAV4qhe5D1BikLK7
cKVfG5FqvehjWQzB73HpdO20uT6BqSs7Voy2Cl/DF8RL/C1bQU8m5soJVMmPfsHIFvXzXm3HwcX3
uwWA02Cg+F4GRncHCD1mCDLfhSckZKjM70Q/ETWwJlCqrpQ3XxIYw+6zGC6vma4yfn13gDUBNM4i
bzqbgyVxCuZ5VV/3OvwneNBi1g/WCeKKJYfdIvwosFDsWgG4jSJTLuVHeI77IdXpr08ywsW3+IeZ
PgljFCBXptZaY/PJymbj6jdou6QqDIBBy1iNA1RJWVCgv0AuJpPGLqnONr2kld5VTGb7kuWfHTXu
GpAPuuR+S2NjqD/OiV3EHJ4pZ+RCxTj9e47DNu4yukBx05RVvXDCVzZ4Q9z1udTIMzkNNz5gSl0K
ZySKvQv2gLvMqawCzXnQzjG+8Njs0y4MWJHIAlFlICTMft31tSkhafDo6I4v33XvGfjgK/VZ446v
7E+k2KYemvTqBa4Na7qj7wlZqzIgmgbPZqBYiMBgYAxbjg18K0ZUwf1/zzKXbRV8slQCCeDtaeBA
04TKu3sOzKI6S59+MuoPHzsEqU9t1/0HY7rqol47o/bgkorGCztDSkGc04fXPuPsz03PigK+xIWs
K1tqdhU3K+hT7oy//ZLYzLh66CfCqb7Znt8irer6bUqp26lOTdKHwUfXEZq8hCcCJEc9lkkNbiTf
YSLG+qo0AiwWDMw0a7OShm8hthRQAYHb9ExqsA5XaHHmeo03KTKZezGDXC71RmbxVLspfURq96IB
eGkBBmijCULvDsQdvlzrAz0DZLcVK898eSHlLGTI2hqovN8XR2fZxz+oaKURxURWYjEfU2xS+jOV
CN4qmBMV2ItCKSFKuMTpwLeEEIUu+kj0FQXRTHWHs8Vk7dlwkMvXBSh5tk3HuBPlkYYRqldha6a0
qrl3ffAvlRbloKa1J1uCt8YMWvk5/Be0Sdg3KCMFD/4Svpo7CoOJP6Nm5d7iBCmV7OAMhTpkvPIU
J0EZ7pV3KKn3hDE2DcDXN8JYw0k15FwMR1cYM5P3htGwrr1RVdMCd/EvjoNZbIgZ4PfQwPg8yfb7
Hxleq4AAA7g9+WfSseE4AdXSYT2RHD+d4h5q1+n9vPaqwTvTS7MbWWXCdzSpnUCM38RvJNd4JJDc
dgkwARklMUC8FF0uIIavlx5iPUmv6Qml+yXDdAfIjm5Pa5Qde6a970xX2APUIc4ZIlhKJEj1eVRg
Qjswvb4IACbOy29tx80VXrXdZkObQWITLf76k2iXnl+0vKnRYPGLtepzJtaDR9ANAFMNyAL5rg3K
sp6isn6u8eJmzReQe6ytzqaf27s30QRbVK5fblRrkkeRbh4q6fHAZmpzKuo9tX2ihir/tqN2Yum/
yn5AETPMM14+2jdVHR7KZ+uepZGSoTTzMF8lFIh7uUMwUtJ7L3rqR87wvJp2Yn+9Sp00RVf8L7de
6P8F8wB6BqOsGyhTtk7+nqPG+GHBQ85mwqZ6wLoJN1l+Jg53oMdDMIYe8woAF6hWmlIWS+qWmlfj
+Id1l0zHZBb9qYShJLZSm0quhGoaGIHQJHXsE5WhKyzuop3huxg0J+5k8PGdFEbJaT1pXdl08BLy
DyBZQrKxzcH9TXRk8BBzqhK5243GvsIj8CQEw4qpW5jbvLjbdajLDr/Dj0NEnvUtS9l6GxgRpOFx
ppwMkJsKHKLZrPG4BkYWe/C+RfHBeOlecV3TNxUSxzDIKLvWarl86EeONtnu06uYR78XSeSmgctp
JXD3YpFqedVl2LCJc8UW1JZGE0L7Efu1pt1MO41qjjjdAwiN8XqsBK43uqLzyzrOlhhW0eY1V/I/
kIfPPM/rfgsgHeEmzDR+xCV7lYp5hzAJ90BPQray92jOddQL3dXby+UKp6SPoPY3sCKaEcSry/Ns
bZ6ugNAFTxgY6Rs9NUCZ5vRcpNoMk5Hyr7EN69mGwzxIO9/6etfA2DyAuj5HgH93QG4z/4xWcPzm
uTAXALBW3h4aEQRaQOYL/PFKmPwHyvu4GLgAp5fW+SwlzKwB65axVGGMahfErPjFaxBFN6QuZh3X
ylBpeRsv+RBWAdioahM0AXkGjkpHuBuzOKP6Qu1qjGookU/kqHdostE90X7+X3HqNtKHxe1djILU
y/1/t8tGe63KCxBKTm8lTxmmIzkEj4zZDhkstwbAwr8pLrwiKHOjuDnWReh/d98rgshQgo3tVcOj
mwE6L7amH3V7adjfaWKKQpXDrmbgKZofItyM5LK8F54R6RVg7tG+xGUZTDoCpRPerIHMDRIlHWOY
w6PXffbYoa4HgN8KHYN92q4P4BVJFeSBA09YE+ETNs8gXzrF5yBh+7IpAVhUtjpkMdWBi0XIHz5v
kzoTdut5Exf8EOCaGqA0ui5BQ3AnzV4g/YU+u0wE8zLv/2dKfBT220Okd3JYLCUPr2Nkz4xukVr9
rPg5Gydu0oiKUmYxcDHvHF2fnigBjmV7SsrdLoyiL3HsQSD9wSKXqf/vsRDXWKIvllc3Sauufn7T
oaUBMENVU/XuLKXwDZwxq1JfycP+akz5Y8ThXS+o0wXoDOs2+vwB9ER1uWEYA9HWE0P0GIk2QSv2
s0xHkk0tAB+sbqElDS1Ey+lVGXfYbptk6heL2TZURHh7w6LKu5Baegm8ocIcvuDW11JjxiSvLxMl
QiooHS6eUazVNJPlURoGpzyvl6Okj9/qCO6MhDpeLLLrV2e+Va9u1pvvQMyChr3iGGoZwvATrK/p
Gghzz2pmpbSjgFkRhMPhdgvbPhJuLw987UkXzfHtk0dF3h3r/C9uEbAUS2tbbvY+K6xNpUlNtPvW
RD0T05lYhV23qj0U6wC3LxoPCCmzjjueEhrk+ryS/fNK8r7f6VufgF012CK9LVPUWiC1aBBiJa/9
/lnvHKu7SJCaP2JNq/tYoVK6SKXKJZK15rxv1X07g2D3zoI1s44IyV8j7UXFj/Zh/OhtZkH1TV18
52WCjlSlxRkMKNy+0f1jdMXUzG0v/GpDTHhC34Ywz+qSPFXQfntgaJ67nOQotoncPzJ2mgtZkvVh
GybOd3AUsunV39bSVuK4JnrnPHiojgebX+oyUClhixnHsUHaD5TLs9l2GBiEFTk3vI52irCmqhcZ
sRBb04XxVR8ICSQOOPEZ9FkMq5qdV4gZReGcQspRCxcfWPjjfw4MHBXDejhppXc6atT+o7WkKvVA
okUI0uClXOM1UZlbUfP3KvEsJ/v5pJNqdm+WB2tjspNwdgcNcTVikO3R14TZDTgg3QztGu02JEMd
mNmncIw1MNE7lGE67ef1iKfyfcT95bi+HSx5VLMIqaBpvtOkxQ32RzTvas6d+tMjWVYtWIAinprH
Q0jHfGX3UGh99HHU/p30gfCfYtkDA/CsJlwof1Uyy+ps4uh6WtKL+jdVAgSkcsLTA1LEyI+bxxYn
STJqm4Y8O344gKCxyyangiv+UN1FfQQI4pAN8jpPqkkDeETzNdWH6G8VB2GTbD2AjyZ+7VvTiJWD
r7yiR7oX6Xesotl83ZtsUGe7mgXtzC4bVuSXVRo7GTqIW1ukqd7Zx6UZUXSsq/EnHRr/nanoFTnP
b+i2yHiCOxORWnG/K5bSlRc4wCyBY3qM+6i3YtGtMOSwrbpo4f9Frs0DvKLBMRFu+RJbErcZ0xGw
PTwff3hUkd+A/+tEYsRsF5xUNVpGN5xEXB/C3Cov/03nm5yCKsGgsMGYF5iqdku7bbSO5UHhn1jz
7t1/d21vV3XjLoxrERmZNbgHExIvOn3+ZA/tmfcIUJ+IxEZRPPrR9c/r5D0T7rzDFCNwK5G3bzzk
06lyfHWOTibWADD0ysSV1yAkKgCH+UiaSJWVvazd0dbHFEsw7Jkcf/fwudGcXxWzIjo0Dyx8ER1N
RqAeF+Z8NkU1P5xtF5BbTA5FHJZuTVgB2VcOCoheZ9Cn/Y4W4v6HKbyeepl2BnqpNFnU7bRZ9ihM
ejChovj55LMxe7ecO46Lk9M6n/jTMqhU4jE5TXUwAeDHZtVYKqsT6/Z+sSKRhYvAcfQJjvWzr9Zw
0kn8xr7UhgxySbcobwp1KrISTgIh6wJx4nVUPRnD1Kp9XH3/TrHOpTb4ebka07hhkme2koZr1lre
+A/8x755O1ZiCiXeAr1LRkwdc4OG6j/9X6kxN+wQu5j93X8ZT9bQqrAgSB1WJo/qOO/mOa3YCptv
Y3KFiIp8zzcTRDPN4lQ/wsOcXsjjBDbsKtN0/KsQ9n7MXUBVV71fh2d2q13VTrqEJPBeS/bJ8zrl
gVUaGCwDQZcMGQ18ldBoRL9bWDBGgGLUY7wo9xBbwsaNBNmSHh+FaFPX4cuOWrH+R24OLYd04oI/
m7NsObrfz5lOpsI8HOdjf03ZIO0Iddxvfwh1auGV2DEtVlV5sINLUsU7A3hTOPMmBilwZSB3BLOw
K3YVN8xhkqIzXiqb6D1PzPe47if31PILBH+jpVoAcz+XrqqckiB9j2yklVzNDFDu/OR4dFnGO73K
ExANiXdzSnNBd7T9hTHgnv+FlAmWgQfuoih14ndwH13OOVjHGvQvF+tRYfXc5jjSpVTLNYMRRSy8
QIw9FNk2LZrhChIjK1DiGBt/jfBdcvpLeV7//xEA5uUE1ZL+NvMKJRrOA3jykcFCftV36qRcIcRa
dZQ4Jnoz9UPJpLyraysy9vLThP7wwX0nqSw7TDci9plMdGE6abkkoOMh+BIT1gbKc6to8sRNczCu
BRahgkW4UJaethgUV2ujH4nm+3IQrTNZ2XBEijpLUC9Zkt0J+ZOYuOruua+v8FT1j6JNbkfIlxoh
hzWi1ceq9ZLWqntx5vT8Qz60rWOrw27h/tFxczKkfZvHqg36B/O3K4DKT/xa0HQX5G3sVIPWaoSk
NGXYgP88LTuAbXeEXDQd1rynLi92xl/O7JqlshZ3zuj6mqLP6yJUlKLfZLmle5Sw8H7zHKjYG8EB
Vc6arQd4kPv6YjXqRY3DP4XUudOqDpv1xxfcBIoOUPNjdzZqGhekZlV90dqIZ2Nkk+bPO6nH89lY
sEfJXd1cdPoy6Z2NTywgD++uFFnCQqSQi/5ig+kGZv+z/FGwtJumnX333kIFZ3jxqVZY5+twA3lW
xHqLhVhYObOVe4dCDtP0M62W48j7OkCintZgkRbHZ0UWQXUIUua18KKoHmAEQCsaKiLqqTB7Kz+I
jJeJoGFt542aBddZzP08U/SCljGZ84CWDJ0Z/B1Za86kXVXIrPOd+af4ThiUdnt3z5vlQyvr3e/W
dZiUm3IfuYuO/IFFgUxcrR5kZLUj1Z11HGaK9YXSo1yFUSW+xKJz7HXw/ko8b8APpX2gr4VdhvZH
VoKr7HjHUYLE0G/XkmNPPuwizYHwWZUE5gifuSAMeUXAE1+lNJC0VrBlPOhhTXeB32UyaP791hG/
JmkNofNKVt/pZ0bSW1efHzH6qYtjdn3dHWqlpP+TNhT5SD3U/SH9PpTn4UNfE1WP+tv4vVBlBREX
za3ZsaEqgbkA6Ts6w/PTQQAubyk0v7euxAYU/Q0PqQkNFqZM21+UlzAr7PzQmqDNRdj8Amykf+uN
Gu06E48pb/yfrnkQJP+t1hvaJBPLc0ivvyPmlB7L8rjsMhyi48DcXYffcor86tiR49qQ1saV8wh4
9X16tz7XOcIsaxF4eP0WP9NQvsDTN49OJOV+Q3Bdoaq/jLlPjguASdb2OuDfLRPTF+vp7jNGWN5x
LyBhPkyixRCNRPlfl+1aOYLbGonCuORgTo1IZunXZpUJ5oTw8vghthh9mk3pCeMq5lo4fJryAQnM
X/Rba/HYRI4S9OpXSjRlVMiwHLcfz/g0UhBFamRFS8Fyp2ItheP2Wmx0vsNbccEkVQW/KWU6sq0E
9RX2P8Xn5UUYWy5CRRTQh9vdyxOsK/hY3lDUjR8qLLPh2X2WeNjfQoC70EAz079FrRzej9sUO1pG
9QtRv1tqGPQYLT+81Jx2Uul60teNyy71tpbOcsZZUa6qlhW79cVGMuHa/cG7+Ipp/p9kC6Lt2awn
GzmIgGlyUp1ScU3u5Up/GZBV7nMoq31qONq0BZSxzwYHnf48qQFU5qtnqEe+Wqt4vqhsMOBV5WeI
MCsPhRLcuA+ZXrDx8PuQyJnWsZXX/XcNp5GRzJef0hZ4OdMiVKv26Tbcb9WwjItwrbq1KoK7WDLV
cCsRu7CQpo6xxSj54Do+1PMvPjc8+98PlqHkWh3rp4FZckgkf3fIlDEcNg69RMFkGS6mZMOsjEOJ
b0vAnQeHZVFOkjjIZS1BkJlOPQP6l4nLY8KnXIY4wyxU3ISCtv7GatRN0mjOaNaJVbzK40bLUVEb
7O2L2RuGlvY9dMHutz23KZGN7rJwBZb6DYSfsCbwxLM4ULNf+z78nAUapdngMh7D5J5SMSta0t2t
OIhaiXDu97lG3bn+QsNITmKKD7qxAOg3odyerxLQ7ZxnZiz06MerhRi+xO5qWWI1XrYV6LjJUvxq
HjIQ4ngIkYh+on9CuomnLjcbqbsV8AG4kD+GOHLlqhtUzc4jxQNiiU4OAxkVOqbqQcxY35cpMhxO
3ScYaU/uOgXoglQ+Y03eK8Lf6CJ7yMjQPL3NRwq37B9YxDtJj02nAzFtBC50VPkfUoBklXNO4k89
hkXiQHLgHajMDc+mQAkq6kly6A/k29NBI4Bb33A0967cH+wLCzjY7fFHcajkhEIe7c8L9OvEhvOa
kGDVWez0Yj3bqEH0qkbTVGahP5y99tJhEzgkylqywGJQc0WYD1ztpjDfpOXdEa7ePh5J2nTytOY1
h4RogLaCmxqy6catvTTe5ANZ+BmCSa4NqTzA37Y47Vbki1Z/MXHs8aXGtJ49onknwPiR/UPTWT3G
ga6ztQ9Jbm+LGFJ8zJwWpfn3jpR/GpFcH+cg7GGevpzYIKYF4Ko/5sUDBQ21mkITJvvquGye0SLQ
IFjQDLoMDXueaEU52KqhP3wKjBQd81pxgNfoxzpDgAGXoz4xrxZ6NtNZFpW/hIWQhfU5VOOD/BYr
RVi1oYPt1Sm4MCB4q9CL4sZg6I/efViNk9PbbyielKRWp9W5aa/kGXOjmfVK2AmSTnRRvJbHv5jL
kclPjjMlArF6v+0ESCeXpsOS0uIUutLcCZ/Cl3k1ikB7j9IXGo/hQgw1yBChPe86+c1SlWzHipPs
C9+qaoQBD8Q/T0xUJg/3FiRJg4192+CQjvJq5/EBI8cxnzF49dP3lsoiqupV4wvVTO7Eyvx01k+Q
Bicu+BF1QQzxoYtjjev3a2oUkngaQIJfianTSWO3JiaPk/4uOLWN5afOFGT1K6dg2mqomDRTl0Uc
/xkE/vdrFqSl4VfySrzTvowoe39e2iVFmEkRi3/ik28qVi/UTCAhsqdvtykJk35iUY+N4nMwCd7u
cDWkdqoTvsjwhmhq+iRoRzo4q6EJrVtXu3a+BfPhdpj8zFzo6OfugcTU65E+2+iGGLZNbsMs0Vir
AQgzGrht/nturTSEJyRrMKuicd6yNLLAjHuwKLRk7otjQaBJM7SxExtn05kF0fe41yLb+Al6Vrii
ZyfsmIaz0x8IPcpDRRmWTbU/lR/gilkTrAxKDbz7Jjc/ERslPYgvo4HmP0KtwB1rgPWobJ0GVdGQ
ftXe7plnhhs+wnlhER71kifPwSlmI6h5pOnr81RsKY2H1gANP3pwmhyOMQL2BpWT8QSvxKkJDJP2
2LHQ9DMtSN3UGI9Px75Agcd/rSUmPHoXF1uaOcF8hNTtSsarVjHP7FDJYtaj368Wvwhk6ksf93P7
kgCMtWiry0csmC/HA6mbotq8r04cOMJRstWW8ehp6Nes/Vy3QbsmnK99w2ndtLKfhFx+8tj/3+Y1
kFvTokBf0bNHlU7c1XiHTigfjf+UiW89l9w24EGXE8DldSJcgcE+WwBTMQlCDP1n/dITWPwjrC3o
asEnoWmEZZty9i2ViPyzU3qIcOa01/11LCyMBMIeyn/2I5pw5owtTNSgG/IhxaNSX2QkYWOM3CBb
O3MevBQ45tKV0/JIbSq54qEI7FoD3wWA3qjoeZeQMDYxYjP8yDu2aI+xxES5ApKa9581TdRxCQ0v
70T9GO/cGJkHK2NwXK2k3V8BCdQEYhZV2kQFgpapoKGEEbSXHOdKFTtMKV8CRBba/9TOUyIsGU83
H5/2Ldspquv3L2r/0XbXArXrHJ1mFnDpOe7Ko3ZDiiKokHIFqbC504ScBw+AnsQPBRccwNiRm7jn
0wEdW2DwAuWL1c/ma8VxHrB4cvAPejOZYpwycr8582V3roliPhuoxf9gG24PL45Abdb5nU4xZ8MC
aX60dR9r6rGhd4yEt3fedG1QuAuJZQHnXpWlMM5v3P2HQHNiJm+LfiDBUC3Bh2pqqp/EVM0vMkBc
IH4ADQaxPQzR3gjGPCQONcD7nW3N+QMU5g6Dqjx/JP94emodCOtEB7dykQYkuAlUCL4vJv2kSYCN
GdZFx8y/IF6huYTWDVGvJ5XaP9kM28r5aYQ7Y/nsZApsLkvQgizDs0ZJWooVmLY8tgoHXOUAlLPy
1iPIK1mMFibHmaZwBo5wMPP1FRrHyyx8HJSgl6F0Uoh8z/U/TeMgiw1ZqNNhQrmYW8bWsxmGSjHp
9J22eTlOMpy7maVVUElDi4gr1tTcYtZABb86D1XVZ+D7zyrZpO9kzfaRZkUR5of0wIQynefZTKcq
E5xA3cNRiSZdVhNMpIql3C3pR7fl0wJHn9mZN3+ft0C2v+R5KllXagWGlaoTj+7RmFK6NNVpBgzY
qDtFJ5zr//685CW1mXqdsZeLGMr1xWAoiUCjN0W7Epkrz+KNDCpWHPid+F4m562oP5kWhG+15pl+
O832r5Oy3WtwYQ3/D42LGQF0ycQ77eYfE+Prq+ZT3r/CAqxjp9wuDDqcFlv76TwJ4QcNDGbDBuVP
Fs1P4Yxu0QLMvQgOr53yN7ad0gwh6bpUdGE38VRul5CT152VhBFtJlms4U0CqCuEA9cE3e+FLQGD
sdyBlyOjBrp8Mdgg823j60RZ7NFHePpzrH+64ffxNZTryPGVu60S4OY7l0iOz7TvBDEezW7s00+q
cnIJs6BJx4k2oi3dFVUgF607HdBewYikZnzdygLqoQzNVnThMlvjcv4EyU+4yAMuWtbQt4z4yuPN
sbh4ts4loot8hcmig/HHDsAcI3Y2rq/PbO8x9bjZVEJ8RTygLmVcUgsjb/X+n3zDu2YCGlsyP405
KZhB+dWDNmTsr7XdiZPxZfjT4PK1tBpz49mk/oJcl5R/BaWEq4ae7QrjSNiD8IEJPh5hHFE5UmVW
FKx70++qTI1hp/2fxwi6XTWeWhjEeOz1a1+aWxHKbhvCdFkXs9dkY8MgswsO6pKOfTaUShkIEPJh
xdxTxwa345lFsd/M8BSEhPnwCShJvV2+RTdNpRY2TPuO3WbAToSCx9w7IbLj3IljPL31JB3HYoPg
54JrVvWAnZOWtDH55xzLBxjWHDNCl3iQNBflDWjYva8/MQsSXkg392b28IG5eopfRXOUfGSZSmHP
rOByepaEgHSNfsiNRTQlgsPABkEGQ2g/+wvp6554Lwz2UM7MxjiFf95aid7zv1EkCBmzcp01Cdqt
8uZtTK87iAFNx8UsfUwVJ4Bl7CoFwIsdje1iR+urJQFZDimUIZ17/nk1fQdCnmbANmHuea/8vBQg
VFkkkeztypXHeeyu7SQ8iM8A1fr7SBgBlHcRkrr7nWJ4EPfRhrYNtr9JOQA0tHJBHQeDvpQ4y9mI
fOZ7CTE3QuLSlB5Bag+Kv46RM+6xiwZg2qZkJKbL4YV5mTM/L4NM9dsL6feJuBUF1N4NmTri4etx
keikDJIuR9w2uZemaMKRg7WrPLKZeyQ0FPsB2FlBIl7ajqsBXVz3v2/dEvKghG9Y9igxpqzM+d1J
a+/dpWz+QdCvBQ/Fx8K2Z/W196x+KG6LXXg7HiYApG2td1y83V7A64iziSDSLFNLL9UTWCTR4qC7
Tpi0ZewdjmvVn1rX2gm5z8npxghm+jvCCeJ2fbWhlcEKKwlR3N2jqsaQIWk8ClXA3m5aUoD+ZJqX
zvjzfdo9f9626lyQoUS+0buqPkl+LwyTSo08yKnud3zMSkEnbmal7NRSGLfCv0g0ywgILkiir836
WBmH5X/sHoXe4ZIvwerOkM0kF38NToUmeZzjchJFTRqZmmXKH+ZAU8zaI3sFHTuLBb798yE/OikG
VwIo1eR6Lq3Pv7g2KYIZUElIjKpsfTFoADP2Fjxu/psyJMX+JLxGyUEQtmOrS2jaXwAt6BmfAEkc
sanScYYlkUENj9zahAiTqtq3GdtZtr1o5Eoa9kzhYBCvjzzk2cJb1LW5zS83UKOUTtRYzaogIiOO
duVSn+4IC6lTt4NA9zCrf+JPWoOsjBXbpRrx6AxVo3l9QJyhoktu7OfTYXQiTSzN8hXUkk/rPcGi
Jmss2luVL+3592bHyhUycXEMtyU9dy3TqjqNvABlX3VPpmeaTXHCfnKnakvVBEVNZLucuufYwZYQ
vj1UXqhiyrRO3kY9V6L0Bf9RJ7ZufowRtVBi1VrA7q1cOO99c3i0gTPBgR49ZvHFXkTTuHhvj/J0
6dze4ml9BGHJ+zg3a0gg1Zi96RklyiDzn46DQcDmfbDLo4R979RCMn8nJlMqYoZyH9YHhKKy8oEY
Q3PSDPAY/ymCs7bMx4J9s1WMkEmTInprSYkrIiH+ukllXR1MvMRHXMgde/vSCU+96K2+BJzcavZV
geYyskJlE8h7duQNXzzwYBK9ONTTz32HxkPiZd8wn9SDham41ic/5HtU509uF/pzfuyn5Doy9RMi
eb9MNaawmbONN9O1f5UyHBaYq7ujArdf9Ypt5tx56d2jOURCl1UreHygTesLoaoxZ3Ka+G0fGeAW
W9UDKWcJrJ+E4dqJvnfw1xVb0hM5mmfuEgg9bcmShPk9YyeZIzGo8hJIIR6q9GmuZqK6Oka99pmM
cGwsmjKXUtc8SY0u4+bCIGGgWpfXe117Jcy38WOlC9w2ZEasvx14RDVKXYi9NUiGSPrbSrK1axlq
oH8s29DltZLAoreNy/ksLaR5Y0izGKOG2CuOIn0v999c0gTDoHt1TfBpt76vwRXIUeHo6WdXnXiL
WRjFzDWkT8HY6F+Avh2ygQAy5Pf7Q/lri055oJUqH18Kbb2KvF/qvrDA8QeiHEVrfG+Ut6exDmZc
LSu32+sYoOqVY9QXbPvzdijUQi6qctN8xZIxS+RI7uE6q7KovQVxLexW3a8sxjtP3dHkZdMnj+TA
68sgH6AfZHLN+rNKo1qrx4145QghnJD8wHB5nyAEhNXqxmBbUYKKDwNmB7NSGmnLSWoUxOhqWtLw
UsZwapYF3EE7YomTLa542Ftt8NW/ILkty9+MJLMDIQqIts/XYKmtg7yzmQJ07TMpEs+sjDLkwUwl
DbGJpRGmXd/xWOizeOAGr4CouZ2WlKqPQFAJHMdtnTx+knSvBPUHD/p1vbuVK8/WzEx1Aip7k+HK
T6Tc9itve+W5g1Z5cRZ1fR93NoNdLDiQJs2iY1Qr+tHYvmFOQdEqfClE+mhCEpSwYYd3QDt6xwaM
Nd7K72uJdO/S8HpHts1KpTCWRSX2hRIqMQaE8oZbHTj4WeajhbQ4yfurPEu7/yP3skuNt4ON/XOd
8sieFsQ8/Rd8NjM9gVaHwppz0r2HZASktSEMrOF/A0/yrEj/JrUzg+qcs8EccaWkleq7ErPY5xHZ
BhRHA/j0Hi93Rt3zylm1mKI0DlWyu0JsTq9AbM1OjeO/WflmmXGKIYqEf6U+YxFiumzsmA/vfBg3
cdrdQOSdjqWjSZJMx2OTSDIbfURuIUC/HclKxQgFuL1BQnSseKROOsixaBeaau8yM1mMSPPeCfxD
AxA/O7Q1Z129NyZV3C710ofJaSDCYgRH/pZf9rhNEwCeMl0zpIFGwrNj+z+o2tITdHfIbMaN6S3f
yEWI4+C7FNGY8RzQwrjYKKHjeasKUSQk5fHnUZIBq8cCbLMlyiCQrG31GPhyheqmRXfMCcNagmr8
/TMjZSFL00tAcL2rKCLd5v5HnWe2hlLe2x1j/QLlyv7qQwvd7wFgGp6GtU8iqXr1HHXYFZfVF+ss
vPVcGTrza12lbuDzJPy7Sz9kM0W4TLOYhM8M2Ajv9TV1qS6R6Q0gw/ip/GR7XYYZhJWaBVLBUr2V
3YUQizE7ZM+z/WqObQaZN8+NQ7IqfBf5QMTVNDKPgmk71TFhjgKtZoQl6+h2MOpO7tMGxttf43W2
4oeL8KwjlkBlOerZF+bZP2xXUmfVdr/WIadQGCChZy34JZ9AQfFANRPjTNIPciCmfvfNraQdfnCw
40opKHc/M+vAsP20V6yLvfHu8EIPIkg9K5U8/94PjyZlU5M6d+/odZFJIjDFRdLH3O4kpZyZOUEN
mulEM0H9H9QtVrvAW4UhEIWc98ASMb05IV51WX3084g1xKlP41B9wxN9vQ3fz4ku8ZN/FcBGZ/9S
IjgHi+sFMhe+9LuuC8rWZ9xbOPHPM8m9ZZzx1O49cPPVDkLSsJTMAJOy0VwhG8s7nOzI39jh73rj
hIjXiBjytAt9t3SQdkgT7crxOnWRxVTvQRsJqinRC7cMX8OXrhU/3cdG2ToC6IiiOi8melkV+fO2
5NiywACyTH7G+2AzA4nGKUkF3d9lJ+GcDRYwXanrV3EUJMGLo+Ez1BGaQNMCy034vTyUCL+b/gB+
D9NMClRJ0L0Dv3ERNaCv+4sDZ9SqfhoCOPWwuZFtFbe04yWXFRa44xSHb8nuYHMdf9ygWzAGdFWE
aY31emqc2jRlYZEnf5FvXTRzkK46V+knWVnhgQotlzHv3eyxjxLdS0a+oA6uB4b2yDPa1CqjWHkb
i4JoMY+dHlneHjIfo/o/qteCLbZdxUZVVVttMw+M5r14s3yCIN/WZh4fdmhOst79Xe9KvrhO+vmb
9uMVMC6EKgRBD2iON+tMGQMepu0BV48Y8UOqjrz9MxSAHDysVQctYFQZQRMXvqtLYhYqmk6qIAMu
9hOYyMLEmZisbPr8CEZ1Y9xhzObSLm5PBz4YVo6S2TnS2C8Do8MK3WCmr4ahf67Gm7ivQiRjjIrT
gCSnvT3kC6tGb38UYjiuWzuIpH56qbF6KmzFNb+xyJ3quo3yu5dV6RYgEggsdGlLMrFD8++LHOgq
iBvXnd3EmQfN+CqjgNnbX+PjzwsLQVDzOniayfPPhXc0EHcMRPEHLUPi9w7fh7uFJi5eCOco7DKD
b5V2O7ZwfeHY4dC6+9TZKBPbSjid9PelSqlsaDiAtUp/MF3+zCXWDlawdX+nWI6fSJ1kgrY1306C
IZ6ZgdslySW5QfLQjFdUVjMlFkIEkw8zBa8NSzNdiYKW0MrNQhX/s63ge/o3LzSYDJLDTY+qhY4D
OHRA0/Qi4kkltAB/HLfOpf4tqsRsnOicMRy/ojVM35m0/8+OA6lPtNgYcxCO/JiE7kiQKrCYP5mk
uTXv000ruNpSlqXJ2ws6WyK3FOMTHjdmHoQ9NEkc4dcB6JTeyD3mHCFjYeTqEYcnCTyys9p1gvVw
DRONDPcBA8BIkWa3GFxWP/oXd3qBIsnymttYRJz7F4pOIxiJqeFTkQqo0btLIKaRDC3jrrqNxqik
Z/IpNiFbCvHJs9oaU6kQS/sPvLehzFlXlsqI0qz08n1frxA+Qs+EkIkBNvokBg54VCGc+q/Bskvn
FDHtVkw9ls8uxUs8rqgEC705AL8jL1kegQ1jbVqWWHeL8nzKZYt5ekgCWUtAukJGCGCK9rUCIUF9
m4jih2AsW50zVV4g3quQzAlsBnYkshIsfJXPECsPDCmJjUmzEn25CBqhSxlgJWQH+QWIFTzduapo
ibhVCsQEmQrEYrd9R0Ef2bASVB+RqJAx6lVXVtEgloULUMDbnOlBKq2R4ndt438a7T0zb2WRMcnS
bG8Rl7O0Z73l5Hm29FdwWXbSd050nYwlVbRvQtfWP7hFGu7PM35W1+NzDdD4eYmB9ULrvKmffVQ2
QzLuXSewa07OZ4huMgBgfNltY/i2Gxx9NMz5uqQ6npfSvaMNjYuByUvJXqLfie9yJa3tsdrF6W8X
HAhouIB4C9DL1Qyi7GrwjX1ms/Ug21buQUTs0y59vU6XqQ1mwzWvhBI+vVCOJSovk8objB785GE5
fA7WqE5PWCO545VuHNEPhdIM/V2kNDGEaoYs99T+0uroaj5TdrgOriMDxlsJp9xvofSM/u46hajJ
ofQN6Y2J6WzMkgFYER+KuTPqlo0iNqG3yS4yFUliNXymtezISEk80RJL6rn1wibuffuGCUPwcHmZ
E9SmoH4+falSOVhngrKmjWhGP0X1lZlqCPFAoXUQ+KgQG7rPc6xFZeU/QReWbCn4TZNynxLa87l2
inhzjFa+rTqdLQjf9ngmP/fHo6BdmmPfdm2UY1fUd1rGwrWzJZAJ49x3pPW34QnmWzSNJl+7cUsV
bZoDUmZR7hjGoid9+NsMvDCq/3qM4xCEqBk0r6YR3a/6AaXeXEmAj4bJofpn6gOIGZZJ19aASHH0
OkTcEQZQGvvU2KIh+7vJ9Rbmn7rs83snvbVu5cw6htlF/nl72V1LdCEiS38REUzLQt+n9r3rANSL
Yx3IzKsZ3TbLKM3BTe0yypTfZadP5xgu06Bx6zu3hem5Uz/VlI4iGXfAD4jXEu51SR3feQ+4KZEb
XkuXe4RQU4HREhxe8B7SfKkXlQoZE+0t/0VtnBUF3uZ1nuqJoZZQ8wu8tDYYjIHAnrpnlRlAoJmT
Gq2i5sBp0bZ7tzDB69Dcumb65mifcJwVh8GggYqHnL/b5oM8pyqn8AY2/2FhuM7TpGCIpFG0WgRw
KIVrX+R94IRZLemq/QdfvKOdw7PfiD3/znGVrjkGEjr1ds52nps5yj6ncFbU7UuZdWOmFCYR7dmB
GpXni7HzFChqM+w5HZMEJfOg938cUMHLPg4Qf5Y8IHkM6pv6RVv/xd12DevgzPdJqKh/1+8hcKDs
n9/SSqVdEk5BwJfBJKOFnRMsIGvsHt1QPEPkziAVjE5GqS4bcNTeTOxz4q0CQzAsFbCFThuJ61ht
z939uwHYwwVq4u9IDOItpZtZSvu1GMlLw8sxCA3twUI/lHAXwtYftT1zeEk0tjVaR+c1aGo2Q+mB
xTUmGIKKqvVvfwef0pWejpygU5FA9YSIrJc6cWMhua8YBb67ZPQd+yBQRzflCD9vRqzXZWo4MXvR
eYQRnoeo4/PCvXHgxqCNDybonWsg6emM4/qqXsJdC5oczaWZyznFfS7ykXNBRT3OFk8l0+SEyn//
+wqZLIX8XgoZGb0pQ0RV0YB1fYjyYsSyO+GsSg+LpeBhUe/jtLzR7y3Xa8E5haO9uL76diLsExlJ
fdtpYz8F/oeUB0FEmPQUpHICQvaTO+wAQHal3W6Klzh5m27YDLNbyBLpaxilEt+VSDahIVw+1rg+
QxoxtaHQPXQKy8cZUVUd9n6cemgMcQM2cExCKTMmbUqHcOkHr9b84MWt/2a5f1VbJGVnlcINbwou
/roZ9KO9qAPIDXAFo3CYzw2dWjV1WrmC0l8E29jyiXc7Rv2t+tUkbydyy0vmYi4/I90cQ/lYOVHo
nuK1difM9WCe37wGSC0vPU6j8wb9NgJQC9+vl/63L6TvONtgPNQSVX8PTNe0ayPz5mbKIpPF9j+j
C8e7j5Mtyf2hKE2FCI10/xKC26mtelBJBdWwqN4agXaL1ExQr9+SRue9BSO90abv25u7wiAZ44uY
klkfEP4w9KgQYq2lPp53Ut6F8ERkVW4u+TKBIcbILMOW1u4aAohecjO/5llhKmnAbnCTAL4GLsr+
Oofu/cRhUP8rt7a+Tioi7nsy8jOKZnJi/7OPKQ6HuvyAIqjFa6OU8+MM0y1bImyS88HvaCJzD4Fm
c4rXD8xAJxS7J3Omjbe4d6+viFOzUHxoZ4fOjGnw1IGjP2cKnPPIWu2iJsdgAxZ6Tei3TSk9hjX8
rDy/nWj7782rApOry1gxKpVRYPZY6o6DTkXXeZzJwAuFLSIDWPLpXOLnmv+AF0AV51uEozGMDO9w
RkM2389e2e3rwAwDB5ea390aGTdtqB0ijoUWfSyAsoJWi9TBsDKx4PneBYf0qy7ZuP8fjcP7JuvI
1zHOJis1twoVaU1oNy3kLiExX4Wm8gvIsRQL+zA92iICpxHoKxQqrgl5hl7NVSrMUP/+MAs9bf0N
4dOkbRFQ6AANMXzCXlDF7HygL/OiChamrd5gTKKGu/fNsidErlN1YJnzwjHtpMWqqqOGCY2/kxbL
9Dzi9itxgJvBY3UjMvi42bo0MaDqbSrdIpr6gTidQC2fv2yJh6I25yqxt7FAAd7gkZpCKb6iUv3j
bxLibKtX5X1d7VUXTGoJ9oow6iQzCbJNIhmwRCRjAhA/tNala+2G25Ilr1KBsUt41utlbDpe30wj
aFY+CKw30Mx7P82NgWKa/5VmEneSJMGOwpO2AtBP+o0ucwbKgVcU0ZG1lXJRArkD/cMTBjeOS4I/
1tO2npnPsN9zmFp1mFfqC+tIfrp/5GtkKo8Q/UjQAvJuBBuOs5KyQN42u1QxaKMrtqkHiJbsrykH
ralkA8hDpdJDrVNHSiiL5MjL1wPOGYaQEJqlNcCYRctBZzNapszQAmYxog4YOzjYx87BZp5/iBaB
H6/1S9slrzkMegS1mtyDP11Qwb9uGgiHe+g5cQuw1j/oR28QCpvoZ98koJ4u525D1NutAs4HqT5p
v/Ya0Nl2jgr5zV6mqaxd9lO9bFRNU90srffvtU0WOHwRreRUWS8LJ4E+WzqHo7SPUhScxyQyTvH6
BD3cZaVJL3dM9L6NpX8LDYUzQto2Fk8r07DTSwpHshyywLb5nMIfM/TDW5+cJ/TuZd59fogfQuse
ZLBU7ztttElid+gY5PmqDZj/8B+Z8gACFABY3Z9PcWEfBY3ITz1BDQFM7BA9RcJhfzGpKQOF7aZg
fbNsqQZ/AFnd3cjp1cEqE5qM/QSVPb8ryoJZ16Vpa5ysCsJQBC4b0sLUYFQI1AwOhMMN+FrRu3Vj
4tzosKeVqQHvITVC9OkJbVXzCTz5at1DotWDNptpo57yIm+rzdZcbLRv/RAhdUgUd+DbJx8xmGLf
PMu6FougGxgqWNg8waVTmIuyl5qAQxQqIiIWbqSaSdTZJvxTBF3k6O8g2Z8TCq9F74nNgCiMtmQH
6CQ7O6xZ2Ww9uD7Nl14ImXElup76Lm8gyxD4ZXcnhvdrcVI0KZ3GJ6HeHhBv7b+9g1tPqDoRADGs
YCQtq4Q7wiIGYAx/+I4emPsuo/gtyvMFK4RkPhmHo3O/gsYlXDTBofbIfdn41NIHJGCQu0QPLE3S
C3Rq7Ok+MuHoATiLiIFaNCBbQWoeHjRRyqVFvTw39uzWxhqgw8KaRJikY83wwhdtmSnnowlwCNVN
Gv20UjWHZIYx/sveyPA2wifSxffKd6S9j669ud6Csj2zRiqSv9WfBLRLQ8SZZgw2wRWtBD70lNkC
Xg5G7TYC4iXjBbQNXmfhPK9tQVimzBlh3VMhrBOS3jAoth5WU2UoK8/z/JfoM6Bl6rlz1p9oRq+h
U9v+nZgVJipBSfMtAfsU6RTfJTxh+gpTXWdJtwSOadux6pe3t870M8mZQ8JzK71tg1mlHSKAMbUi
HQpJhAyCrsncuY8jo0db3irQX+EmawtmUg6GlLDQh+6Tr907hpbVDNBGTCWQel+7vkTUT4QUCrBh
neZeOnFaWdj1t04B0c2uahY2qrHonyJwiBsHOU5V1JhAR/zCou3s91ZBuAY/oC7WwKDBqdmIDfWX
rNF+h/OBR2xIc5/BLyVRpMn/c0S03lV8HOoKURQwgat1KDp2S6NsyNUbM2V7UhgAduTAtndeZdix
J6Xt+mejm8MDgVRGxiYJ2THQmTnGsr2dqV6fAvjc9yGDmUA5kUxQlSCd+/5XjECVgVTrum2Guw8x
eP7+m3kOiFEIsCBZtg3FIdP5hJh6ej81ExO7sRTXB34KCE/DGGpnV+tjIJyzuXgW3ZOA4I70RxEd
pUkuZTgBVpfPOafaVx0BOBn1QnRBuoEhOPPnbD5I7e7szSwZFfQFKaDRl3JpOLHW
`pragma protect end_protected
