// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.1sp1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
OaldPId0uu56p0JfFNQslnD+YBxxWHWwgmGMVfjf4h67mlISzSkylytw33gQzhbE
sviMA+CR+qgL5IEwNnisNsmX6fu7b6L4MCd4xx2TW2XTtgC8KQTR5HciQta3RKKj
5vHmGVE/8Sb/AbwN779rAbdcAj5FyIckEEKUyGFfnwEQlvOeFpdGhw==
//pragma protect end_key_block
//pragma protect digest_block
FucguuWOXJ9f5jAwSNKGEQNjIoU=
//pragma protect end_digest_block
//pragma protect data_block
0XZeIcifyOK397kbBWnol88EYvaSf5D9R8Tnx/Ydx6+0ArrR/WTZTuPUKCMyorZl
av6P7J97Xt/wLH9/Kl1OL1Axm697uAyEXhctTnW3BmXiM5snKX0voWprgPMJVqIB
O2HJH4xlyUjpGT5qcbixLeqhxsFb+NMkyk+okVaCCipOVht0CLvA3assLIVo0JsM
x18KQJxId8mAOhpcCZi56QPR8xGM1Hc6LxYqRgZDEAhh8cOaBHfYW1v9BA2j/Tsk
cry4UGOMLeBxs4STbciw7TkJK2mMt4QjBJhArqwaG04S0E259sWuwDLtwmnGlo84
KyO7qkRqnIYOXizWxdP4kF6Y4Ia78MzwKmUBxc//q/9AXdkBkEmt66+fUAfd62pl
67SI+qNEpK1M2y5lmRM1zH3VZ7GpT6TPUUx2SWDXkOsgLv62zdTHHSK158689U8v
bcXZdVZS3SvOVxylOl6ZIATivwawGTNeRL3O9KQg8mUmdiosOYfyDngm5h8DLjwg
IxDvfpQnU3YCNmQTCjHXV/OC861zH3O3MlttY1VdYAmUDQaCAn7HmY/J7GV9s5Xm
ofv17e7bgUVPMnrOMT6ZKk8HXskJ9rAUW2KDDH6mFMPzmW7KFBnL4N6+ISPiP/EZ
AXZme5tLbVrney1Y4NviONUDO/PWYy7Nx93o1pjkFC8tMMd4afClUGzTzEBIIqiS
Ua1EuyXqQ/wLCOYbRcyn11kVjXBfQ2QVjXmNruvs0AsKq6skAsgY9sn0HoGpjqBf
kPFLc7ISsAF45Zt5/+D9QV2MdrxnXtDe5y70CYVgU4qnKwbxh2PtqR/1hFZcwlDU
0srM9DanlG4GyW4HlystdCz1BzET8MEDhTrD7oYpGkEywuH5s7nvyrTP89YupQdr
/rOc+d1IK0Ogm462DQykLRMmTLKUPsB6LHVbKFJ1XyxYywqmM8GkNEWfXHA+Hs26
2ECjeffBQ8EzpvA3IxsMvEfbrIgg1hwLuwODc8v7o3ZEV5BuzHGNY3Bg2DFLv/jz
d8k9KgahBx6f6tTo2W/su/1wEgqkDllgV68KbZEGiyrFiGZhFpLU1QHBafHon1sS
op8hIybWqxRidCnA/eAJWR3AzHWsfGsyOT50vRyoBv3Mcj6noHD68XYU4kVVyCd1
JWQqu783pB3hGt6i1rNrrzdjnkidAalYGi+SruUmL0A2slRRcIfPY0XdfNIFa/+l
GZIyPggkNqBzKrq2cjRA5kpgEpyq3Zt1pjlIMMi+P6YwPjc4E23RoSElajPJtnGQ
TX0Ui2OMRmtfX0tUhgtanvToiBykDwyzFIj6wYhokMKi27Gh2aKPGAed4Lvc3rv6
oV9nMnQfNOPFx6r0LvxwwFqhyPrIUDh/JOEK0NYltt4Md5/7Chu6yiDq7WOgVeUY
f3Pk/y5J1bY239zRCLN4LxRvqJHSsG7SsrUtpSRELjO7HFzCOW6D+9Bia3f1wCuK
jJ+DU2saHxT6tUQgYAEDfvWqnwrwe1Et62G1sgMhf5fsZuj6CMoKYYtOfoiSduT9
jpZI1+5vo98UA2VPBEsGkVaDGOvx/7nr5t96gOlL25TwDbHGeLelONcurA/Wj2Fc
uj+nPi2tQO9WMGvyKPiyWmmMol68GA0CH0N5WrtwFtVn/q7SclaB58THySLnxnUu
iswLmeWN4tscfMdeOD8qmZC88NBkmxwrCQ5ubaM0TieB0GmNohrqb+m+/QPoV3tX
/bKg+VkAoHXUOjHrVPm070E8r5l3ccWnPfMLi3BeyGANAYYGjgdwoy1n7Q+FT7Kw
+TN8YFNdPwj/I0MJJnWTKA5ebG9v+wdXXnl36Sq8WXmLtt3/msXC7vp7cMs3ck+y
Yqm2NZh+4I/9yCMENJBoC97glkn8yvkvQno2LQn+9BREg7x8aSBLSgyFRFscCUF+
6lXsW94RtXDQt8mRaIsHIEuRZbDDP0edM6qLAug4CFhdmWUscwrVgM7G7wW/5tOQ
b0Ke1fuoVlAn6fQeGi9hNlf5vAIfTxSEZqkFkX/r6eaP0yKslWsPsbzECe9yfdwq
fhGiX+IVdNI2HbtUYwTjS8xD65HIigKhIQ4Gx3rab5+k2xvmNrtQLHs/IGMuXMeF
fy1+D8hz8LRZzMk0fTMkGQzOXOIFFoI0MOS2pYfcVQLxy1eI2hDWcy4oykcg4un4
TAnHKTZcQTX/4+/kj3vzJ/lxGKKtm6GvEpyiEj4ga6RDDG90e+ZcCfg0kDu/jgHE
x0ahIqUD/OPuFBZM1kaE150PrqMmUlb36r4o2LMpCbd411M/8QAbRda0oecg96W9
OJDokW3rYcVOWHil+LrIEHgHiMaZwHnT0gS51Y/QQ+J1WOFQ+Fl57XK1RVb8MNCj
INZeocIvICXlsEuWCvHIlo766zQB1Rq4oXyGxw2kUjIVIE7PkIqsprkqOwkPGr7k
8HUQe2tWwbCoF+71leu4DMeAorNdbqtfsjobK+T+TQRISF8+3hS5vYXtb9TJmUct
BoJA6Cj2BQqtDSJRLrs/CB8ZY6SFds6mbOaB9zh2P8B0wfM7aBhEfTIeH0s+yJ1a
woGzopyT95i4BLAdgVxOZYH7hjhUeS3ifhoHAs09Sp5klG5i2HS0U9qjvUwPan1x
3tO5P+ZRqEujCqdMEFrGVw1SLzKQtbyIvpfyfQ+Q+pogWaxrAzoNuSsGu1gBxxY8
QH5gyApFUtvS9DYyVTxfo+QGpy/qvsY7/CfuGB6av28TOftZ6JhRw8CoJiFPu2bN
BECsUnkYyFyOuZTGcUw21fSCRre3fBF7TSkOLVP+zJxXHYSChSKBZFfhTZWPrbvi
TIHG/VeRvzY1Ph2QY/N6sw6nCjNrnOrgxVvb/iNiiyzF6XOLhYh4aenXd/H0Oa9F
h7pxL6Cb2Ge+Ne+cq5qqjS9sKgC9C5s/n+jz6Z4IDc3ucTE22uDGTTEn2UIRGKQC
5fQeWrfiYFG89ZV10Gl7pOWzPhpuJ9JWuMJf1NJo1tmrV0JbMxE5Mj/zmWwX69nj
cvbyWbznBsDkhhQKWbM5e3uFobYOBYM5hGCKv3KfhpVHDcGLZNb53Pi5005jDo1r
3dBrwwRAMZZ9yGXP1r225/wFQqkb6FM60l+jVTy4uz9mUdRkLtIWfNCL4hzl2dB8
xUlb328IrVOGpWWGanuCr0tMrh5zbojGqPraxYpCaUzdIqs/iTOAvb/fIOpCb3lt
YbCze4LxbNoruCE6QgQLxRkUzeco/0chM5q8AVmVNsVzeAib8/T9d6Vw9st/wSJM
Y+DOFf7QjvfaxkxZBJO0aXU5OKAND0OAGpfDwDbX/OPPCC67enxsvZQQvziS+7p+
zqFoSd/X73D9Ns4ImwY7vMvPF0Pm15ppb3i7mVlECT6MIIMTYZRb1OwmGcd/bLhl
C7MIwZ7ksRmxxoM42OK8u5mm5/YjCbp5HGautk77IAw3s5nw2Y2nXngTjpUvMNmx
/Xtu+QFur9mypqcO5VFS2/Fh6tzFyQai46jJh6UcPI2CgkcAJuoCgbjeJrFVdqFf
5ezrNqDH/2Uh3SiJPq/Lxmdo06Ct9W8bnztMJzha6c+nsGNZkS3jcKSyQWy1cL81
OoyKBrdfg4smt3QZedDfzVjAkbU+fNy3PrNMV0dwIVk2i/99qeiZWDUi56EBeldn
Jo0n8/JWHG0wDKdIjUeIvAaD46VCH0r3n0cMiNKdTPIj+HeXcapjfUGoFyII57Wj
BtnWLDUh1XnkILcq/t/0G/egGNEEgz4H43+M0kQJCWozUw1G/QjXBc/4zDtKSrJZ
fXom6PgISpi0KnbGncKstuUa3v1qLUXQfwjzVOcmk4ip9SoyT9rs6nXhOkjavCaN
5ORD29kEOdv+K/ipaqKnnj42b7IbW3IxlHInTjUKduhuZQkoyJwdCJsX6H5OfnDd
YnmOUbfh38rCgTQxk9qVKDsDmL9VDHTX5B3gRajfrNDFJ/LWZ9oE3SsVt69nMuoM
k3pMeP/+gbMa4ZtHmAdsUKzcu/+0ouciL6cg65qOk0t88cUFEbVd6v+GitGJ/n7i
ylnnjBTUC/NHcBj53GOnzkvJ2DGDYm6FUP47x9W0LOQGmpM6d8EQwbxVKMjSTQLO
I8gSZUIdCd2FgpUTVqT3YQzrib042VWOIgwHcCvjLWZMWr3E/glnGm6pOp4JAboR
OYlpLlu8tRKKksqagnHsjcBpp9N53kXH3PqDZO6IdC7b+y5n5hmSHLK923gCUXMc
9CInBmHKSSvWQBeMmX5zUKCbXJQp8VLAGSusHeCZveeU0m2nd5oMrSsEXXNaR1CR
02VyrPt9aGgMZJh9wI6BWtg540wIGhtm4X8IIIRxx8GFtihQfcZmKT1sge6gynYA
M3VQymw6hwCnZtxwo8Yj4eL8cQuBBEcYPStVT+x0O+fMgrQpc2AZQTT4d/72Inm0
YNIeEWuPQR9yno14M3VH38PcH/uK1eMN6GGI3Kve+usYA52CV0EwmTll3Zm7hk+7
QqLzSDDynolSwUIvuwB/JegGTaTNjOAEXVRJefeQODlb0aDMVk+8Yf/Eo4aeLuNu
g85VWq6lPk53vX1GdtjpYqrxaBCgIQZSPivCNJW0L8QDkcctpUTzMySa5uHU/TEa
8pxIoYv7l9H9Djp9fazwtg+VMKbLAsLB47irPx/UitKpjVGfgPaB0kQAtahJzINy
3ED6yrUfv1STwiYgLiprM1+v8EsP/AWQNxNtwTGkBVy6GIiVfQvGf80Idliz3/o4
duIOPQZn6qQV/7bDokxG9KjoneD4aOL79heH8xO3Io+1huGfOPLlnND/+vpNX/XR
9nGxcuYC/fbDzfxXAna8/JQh2Rf4zwNPyqNp/p+/oE8HE0bV0k6COYGSpf5O5sPt
tH+OR+VTVGfPT6aEluU+VFMuIONpOR0WP09tBRorzhl5tJwejjZbEa13k2k0j+gM
3jnuDgRjcFzeM7zOVR70twkbzrR+T02dd3hUmLDj6THjfPieuuaPkPTTspxlyKdP
JvjKeq7/fWlmt43FnvSAu9jhBGm3s5+umVgOSbUDNk1bi9xE305iKOLJOEUqTm05
Le2YHffH5XLOTp1PNry5ezUrBWD7NcpZiTg4V1Sx/aMB3zUVlykHfVv7XXiVh6Ah
w3whC2ZRaNi4hb9wFZm9YUNYm8Uul3ZAbcn+LrQPN3aH4XSLg11hiBm2YHR9AASq
bQ4dMIbC6Taf0mr6vfm2IYq6wCq4MVp502Zk+73gDxAR8OqSNpD+2lehSORDC5BC
7NNL0o5hdII9Km0x8qtjVd57sk2vAQK+I7fQ4w6tBjRjbwwOPXc3YkeVpP4a2SZt
6q1DLQ1Ph9IKEoQn1KYnoH0aAa6W/BUcyxp1D5ORrbQB1Q7TCJl822pyGsiHrLjL
zzmeQDC3cgoHicARuXi8CXPw++KeqYpiCUppFjVbjyX5QQgcJAQstBDTzfvDjpHM
uRvMVxToQYrzD/NJKwZFbbmh5JiUkSNBCafjXivRRiUkjJ6/r9zhPy2FVjhvu3m/
t9jlmNCfRPs1twQer9QKcfqbgnBWW7wZflUwHN7rUl59qDLlgZEy9mVuGhX3hDwu
M+cX+rAGDmXScCSP1VsOJ6fO8tvjXchUDErjeZMzbuie/Jjvjs0Fc+YXtmFmk0Rv
D385GaQeBo2FNcIrw6KPWHU1sUcJ5qVeOqij/nudgoGj8THKFr4KF+6KfhUsWIwI
3DAbRCkcXMqnnAPr/vpqKS/Ep+qowcIhK4Cs4ipejxag43i7tq9uKMbzdMyniyfP
9/kcUdLN30iZQ2kLNDBtBYsE3TJQYr/C63Ctrsq96Qy4Ak0BPv+UhXL86whuhkBY
klkiYbMIe15nzxw519PRwERwbU1flgufzF13c7QLZ1a1u/btLN0DW3Z+fbItKf0N
+oFYpFN8gCiIV5KZUFp7QETM3u+Vv3d00IqUghy5WUpNebSG7gk9F30NNrMK1dui
/XCsuQdrg6VErio6OaHNrwt2UR8xA1UBTx5HOPrZX5XYp5lsKmzlsjJfTDyQarz5
MWoJVE9KZwHVl72NQc/5QKq72jrY1jvduHkkO9AbNwBo8+puQjJLjm3K7JBkg02t
uyVO6VaDC6YqvHAHZfeBVFdueyDnvmqhxQWaLkeRCoKG5dp2EQ0e+GvP5wyxA1pg
nwQ9ewmqBSP6wiS3C+E/0jmxoGI12b03QnORSJxbIJNkBC3v7AuKXuSld/b/5Tbr
1vUWUCCpTE3BkE/Zd4jS+J/CwyApt4LDIBxX/+3s+TQslsrG7mEV+kL0JByIle+o
ErBvqklv2lYbNOxEGJyemRuHoBsRVG2CwWxtbsSrjRdoNuOXHwcnIQQFdBz1JesC
0Eh70KXA10dnXNEzaAX3adXCKtpyHTdXSUtIQCcL9Uxi/McTxgKFd4i4ifvyth11
YxtuDrD3ml+zWUkp23H3LC3U2VzAjoJ/v0/Z4bNemye2MK4Q4Ew2XI/6b7CzIHcR
tZ/HkTS4qP9H1N+kAn5Deyt8erNhG5U444gvOwUHP+HHrrwDj/Tsx/uLA7ulAxqk
Yezddj4UqtdmYVtEagNRT3DC9ZmtLtsMkgAX9nd0qBJ1JCkifSW/byTsrXsnldwM
Gep5pkfPhraj2WdGStsEXfQ5IHhKymdrVS8b0V3r7JzQAVfqCXWv1B3S90fzH50k
MT1MrfT5Yp7P9v0LH7HLvkl4yVDEPpu2dMigKO6xXwP+koS6ikzOJ4cfOHXuHJd4
nAPr+r+2eujvFpww2i73VRA4P5oRUbssN7F3+JfV1+uGA2QDA6RkrSeEOTzTT78I
XNHuTnZ2VritrVZO+rerhgQhjijsaCXe8ovH9/WkHErd4BoLbajhCOUQnOQuKEyM
t1qhwnJEwXfKpq/82CuSSpgJU+KeSp/X7RDQN9zlDEx+DqjXA8JArGB8G2Hwix1K
RNiqvkI+44SDijBfHFhTBy8XyVQsdEcB/zFhybdVRUycSygutcm/IclbKjx9GZbZ
Az1jTFxWKXZDi1DM8GwYS5gq2uLzaoB8S4rflN7w/u4tIvzCQJWJCmyS2owtAh7t
Sz0u9rdJ5l2UxgxPYdTrizmib8nd9cnavkVj2hqUPfQQzLxct529yWx5/xuCvUWY
eki5fTcZzK1TuW8mE7CLKTw1NWl6DzrIBE1M9O+BnT9Q3JUrRRCNOVbUdyDaX4Hg
BBVy56dN+m/OyM6Py3GBdR+TH44OC6Qtip7bDgoNgs1AZTiITeHzWekoncBXXHXT
8kmln1svI2k/I8NVrBx4zfC9Yqps6XkKLd1cdI6sJKUYfGrVBnbTt15wsHsPtnIZ
o6Ogo5kpuQHlCzIRkha6x/TkyTESbbLvSRUYBB4nV5z/T7s/huB/alA3nFdJSNDo
EI2mQtDk+NfNgWQ1riXv95XIC6RxNNS5oqzid56Zt/oZlxEqaE8u3zUxqVHvCmzZ
/WNfHSC/GqQwqru46SFdiFONbArudgbQ74kgwhqSnSR6UuAZLsNiu8VvzaN6m1AA
9GB7XcBwrYCi92xdvPaOBDFVg7+JjAFR+wEajAi3JLPWMvEyaEP1RpE06tj1/Fj8
+wPpPdfyJYLE0A1wCiBBbUVWfXCEJ+/dgdm0NEjinlUQHEyaKLrQqjQdCWpLUC6g
mGDSYTmJIkRj6UIQ2tOUA+W23ytTEGagYLbCJMpewdUvwZ02mWtiuF/w8bEHct8b
HeePA3JNBILlHYwgbOc4IHU9Q5sHI0Lq7lZPIQ4um6WXmBjB3KM0+RUvKPLHBv9U
evY0LZQjyf+1zaSPHId7mAMHdxJjH8xgfcBRSTzHtp5rLcupbg8sjH1ixfmRwOrS
fD9w2tm2c8WwFJwUXQu7AUxJZF6cVRfDL5+vVvaifTYCjvoFUa08i9t65EwcdLV8
Ck0EzbbVPB3n6GJH0/RnEE25IbigEYENMtliYA3d/cpHo6RUHPLwB0CajB6KbC6t
6dbM2kGK1xZND3r8hGLPR1tk43ptzbi5q7NgABolmsFCbb+5DO/rbNqCZdDKbD5u
jNIyeTDXiXB0mupeHLoN81oQU9ts3lSFjIXWqfHnWJQ8+9PPoypxsp1NsW260rPb
lxUT3AZR4iVeUlJ+bIhgQ9xs1VkPXDmvrK7FYZD0e9yFf3mp6PshjH1O7KyWUXTs
QbqedODZM1VFIaTAEsfQ72LkMy/7c//3lmH5c8wzKAQgsarNjSpPnlKuU0+5utne
j7KJZgBIlkfIg5xrMG4uoDr117qat3HHe2lOUfZwgX1hLX/PAFLlbjjPWmT/byhz
q9qH8W1FrF4BSQG03qQ/KDGBzcMBU/Pnjlilj7k4MxGcmIAbOY5tiHHYltLjR0pP
gAvJeSUcGczkH+cCkBYwaaLX+fD5Sm46jnvJmjUUCkW7f+wEKwNWyObHlr03BjTa
N7TbwqCRycHf84B1U0nl3q3pmLYhvjBOSqISstKOjsTvHVDUNMMnecWSs495oswW
Ua/v2DpVy8LX6+HXlDaWex5usqsJmk+AqKsTpVqd0UoZ+u1JgESEiHcsmDZqBPmG
tvBwfVnn13oqnHBxyWxEnF+IlPv1EsjBsri4KiCI8ngcJLxCEI6hNHn3Nx5sLIsr
7ztNZFFPqA3ov4Hy3VORaW779UD3Shct7J6NpxWxU63LqzJVyLFzYDg/VM7MxYHy
Xr6J5l61BbgkMKWcLd1mcIlEiBP2LvZjrM9w0p/Il2JmkyNk7ik6jZGA9PbKynEa
0n/TuteK86rbTtmmAUEhJXCQeeTdx0v6SFjh7vekrCGdzz+puwAuvxuRtWWB4W2M
unM9ZxnMHlWBPhZCIGaYjB+exhKPZpPHVZeeXGUq+1hqYTq4CQ0zeUdUAc3fydCo
YIroS4NQxnT04o15iVd9uTynd8imxaSnRawXBbDRu3bwafzs4LcaQmRBoO3uM4xd
fKvFsrCSh0XwRWk6pDjIieWK1MFdToeqM7koowDObm95DULAFIzn4hVMVuRrKgmy
a5RNC2ncZguWnIb132pl7v09b0KESJohfNdYeGnhAxqw6mY5qZ5Sv9ifW4qmH/aV
QWtZcSLqwjuPPBWQ2zVjPqFX3ovClhXBFNI7N7urmi5AHr5PEBDs1mxXISmAgkH5
/0hMK9uEvooermB0fQUaUQx4JE8ZnOZ/cAlgJ1M0zBlKiKY45uoHeiv3eHbm/HRC
6fv/DWkk96DJB3NBe4M/sC1ll0Du/ItoqcgUVwL2h6kCDF0TZgjaEntT8HUUfDZy
dqcmapm+aRIDpwuoVMBNp6xSG8JIsftTMHGQW8S1SMQelOxmVaxKcLgLoVlFoGFp
9bEgE/dK7dcL7TxHYskQiNOKfyqDnreet11ERyGLGKPyxKDBE4fu6RtG33aBMxlh
z594ocptzAyau9PXsWc+V3qAfusiNg/oc5VnHtgDZq0pIA67ZWuIVFFA2dsntpVl
j3KB7Qaip2Y6gQqeP/qI0j28tnuNQW2w+sW8rMgbUM1IjLiiqApuRxMmUf8LGrlD
xb+j6L7y1Vjd6Zu2By3QImHqSDVBaq7J9QSWsFIBePy4wOdAWR/2POMu1Y98pqld
0mZ/2khr1X+dLmZ/NlhXKdTOvTtzEnF7lTAbf8FWTpJzNOXIQrE+Xb9xi0rT0RYy
iCzFrbSyzGJYx32ZXe0aZsnotxaucIlIoTEJxvP0yMaMMB1L5fTrHBIgVBDJGMPn
hdEdlo9dwtAAM8jbjM2aMYiN313JKfrYkbFuxwgPELm/C756ch4bvsQ7JM+XSqyG
i0QQodPS5kOX6DOpgXKofskDH1LaLFDTq1GGWUbwQuT1yfjNdScWUATtMQIumJU2
ZnuzHPePKwid6SO37yoLpBk+goxyXilmBA/8d7szO/pCmMvLjFiHc6bm5S3GEb0o
HWoGF4Bilwg9Yyil8q5f+5y50+kOuTeEeK/XSTFdLr31/axdTfVsdpqTwWbqoGkh
6Hw1gAm2+BU6m2I4RoV7mKGG8jcxLci4T16T90fi6JBv9++EZDbHUFVH4PsNZz0i
EFA8/uoXQBVMTgUL7HTIcW6Ygams6RqgdiawR5KZCxxp0+fV0vL/GAoZAnFv3QHL
xwwCd1Ss0h8pOHkrvTMTVwLCiG6v3/YQ+ZAVitHEcKAhSvYomypZfTquIDkJEs6g
fWxFLviZaKS9ZJAkSul5UQX7gshbr1T7IziSnXvUsypp+nh1E+IZdZQ/uQaUSLOj
kMMUjv38AluGgmb6hAGTze2gTDWvK5Jl9MJyrNs5VpEQ+PHhD3E6ZCkUTZTTch54
P5TqZxpSaScK28ROyig0uVfqmQ6vswOmmo4nnONK0JypDnxnl7FPE9G201RTOvX7
obIRQwO03dLXVGmvUtzmk9yOSFKKsCiG/mry0oc7rYvYuBCuhbR1qrLZepgpFsm4
HQsutpT//IvBG5cERG5TrZTwjrwB/HIQGlia5ML1xe8LY7N19TVzxgAZwX4D+9DK
QAsD4o/OJFKfpyc0AkVxaBFtYoclH24ub8Kw8w+ip03THf7q05MhVUichHA9Y+mb
PChKKvxuGGYx+o8127tIG8xKKperK11EWqx65iRVrYkU+NDwQde1IUUsyOEonePV
J2v7z8N6fMosXgasmlPw2a5jU2l2hfvg+3cXWxGuJX6myUKuEJRBvd+E7VnT4oOm
RXJMaEy8t55Pm3w2L4c/VsvvdlzED1Vs4VYa7ljdvPWLT182KZQZW3UMMg/bND/n
V2vjVTkAX0U1P/RUoAontkosflyj+JrmosiYCnvDaYuRo0adp9mIY6JBLaU+VtxN
Ps697+bxxH8/WJLAGzSeWgPnIJrHbpNGcuPZYquHcerH4uSs19xMgvH3vJFY6k8K
rlxXLeuidbBDU8ql7yRZDywZGGwsGBHB3mP4MSgURghq4l8GWRKou+niAKZa8e7x
KS/eqMsTkKzz+Zf6Q4j2OpTd0RTPH8BK21cS1+QjFtgIi4q1s1hps7dwQHqeWn+1
2e03tLMwsyUZ79KPu5RxT0M8gDsRzyGhFx85vLsakXu66E6K0a9Qqs1Q18Au3PHF
qoC2QWgPmmeFnfENVyjTMprLQIpJgVsp9DgouWYyGUC+CfBTmQ78B57UynFB7bST
lB74VGL/8szzmGNyY3OeMXOuomRIzvuz9XO47Ka1DmwlQfBfWfdzhR8sdAVqWC/x
+tpTBLJETJCfZ/eCi+/rTs+Ir7E5jK8hkwNvnftKfps36q1GzaXOdD+4F1t84WE4
iiQ/busxwVg+9DW1qhDw7p+HcBR90D01iQyl08brNNr1dpKvV6zJ4l9erneqft4Q
d2gIUHRz21mYGelekvfjqlpcDysvsRFAdtzAOwJ2ckdHR/kFZvDXPbkPq2GRYP2y
B0q7IV/4RrsEV/YjyqU980o7YkwF67jVW/SoYij+jvnS7xVZxOdpfe0OHCJs8G4H
B1EpB2LpY2H2lw7tIg3091T2f60BvNOu/Sj8SE8kcMyYcf4VS4VRku0dCusMFVIK
3YUg+bquE0/2YCyTEUSTPcj3GRKGw+GjXVURWUaW2QsMgK+sV68pLPkuJ69wYUYR
nfIfF7N/G3SvTkrTAav9zJO8F5e3t8/GUpvobyFxuqcygMMGniKi2ULde08KF3OZ
ZQSJkl4uIl4PNxQyelar1QHhwdoNGTUBSGl3FBRINTmQDf27/UrF2ysX6MZJ+fN8
1+s9ELCyC5X2uuFxXvTJRWpEbAS03cZgX1e+S6UzIu8LlCTAkWYSWQiqg44HVpXk
DuVDsdGr9Y55I2iTHXFItuiyVHNy2omtETTlGlLpDQLKOV7Dvh9jJQHGaUurCXdN
nezmTQQTAefTiLyYcqL6We+KNPNTflnNbYQRaPuw6hYXiiwTWp+9riZSD8UGLNkK
vm1hm8b8qaRLDdstzTqM4xQ5DZP8NJxLumVtZ6s4Sv7TIkHc2r7gwqvrP6f/Je3X
eCNvruWbrD2BbKDyjoHYaCr8XLhZc/4EgmOClw/fIR+kNf1CVH48ZY9ogcRREJqd
N3LMPLHQC/PnTn+JCbRQHiWbXzzQpuOdAGvN0CXyCjmkPj0NI2oBYeOyOB+BTCoO
IL+swWyOhPLRvgbIT6uVkP8j3sHHDLO+C72yCahAWLbAVooZSUewtWRwZpG8+zou
P4sG7oKfs1zId631d8oW91gIY47AScTlzyemBkfBcmN4HeZJi/J+cCqJcrqZMnTO
B8A+EcuWshdt4hdA4PzAXGbM4gCCFBXKHgTGm4rhE8RQP7YngDhrq1aTA9Cp+Jyh
IVD+Zy6wOfykY6nw0PKkMsG3nRDS7O0S6o+/UKr4WrgtLpKBskaty4Ll/6p+MjfM
E9jt3lb1kk8cDANWQg653yOm0Tazy/PvPEtvXli+m5pWn1ecGct+Kfny6zfD6uAW
TCGMt0z6GArsEkLkDoAuz52424hApl7/tpHQPP9Nw3L8xgL8e2fQXDeTFvBE51XZ
Ay0oqTxKxOMY23CIShXUiKhilnAvQGL5sVjVOB9AAwqhIfzuXcSlMAYTbL3+kzXS
GhubNLfhQfVN2DLe/Pk3TLMkXg8X8KaolilBIIHMkuA2P0KDe0CF1Fe1WpwLkMY2
00yfaM8FG4WYFwIS3f28Gsp4ORrS5SAS5WMT1vw9P5ebLRpgrj87e4V1GAiVSoxZ
i/PW+WdoJQM/7Of3v6DR1bBJCYxtVI6C+E3b17nEWA3uyyUFJ3N+HvOVX3vFHsVV
zYR02vc0+vKfX42xLiZ5a0OtsRfmozJIWXNndnZY8ckQJr8WtsZLCy2GdtGSGga9
Qyfwl7igqhXoHuwT0solALLRgNS3mJVc7TYDxMTN+ldTXNrTepz2prOEGImcDvJt
a+xOPVOHT7CsUwjwGxNYfGgkHLsyKpH0+C4+DLsKNNzldGZFIBjPxAiuHxDDpwxg
fTCHDWLY/oTmYlSLd0IDLKd0ZsP9klF1Nd1wpzfOjD/TTstnRHgMq2OfF+buwfSi
HXLiqG5TMted1UUh+IsS6cjDifVSg4+j6/844DFVbCijRX6kWf2QuFefx9cXHClo
l1TcJC8ZH/XHdNB+Aoo4KQbWhV75XrxqA1AmfLCt72gey8A/E6PMCBWXk5CI4HdV
1M5NsZOFbojZZsdPESK+G3jphdik0RIagnihpAI2MhVsFvBRgOtahRXIlSYzECZ0
oDRpDm2rzuKD3LpLTPh7sxEppjkt+6ZSQ+zDzS33BakJ5bTQDlrV9xk1eC2Crdls
TgOKhOq0yWk84DVIfIKskPcOoKgfr+0hgynjvJJbcO6IGh2cBzo/j1OsTCig+ODC
GN7yH4XhSykIv/a/uxBl21spGqeW1wqBFDN6+2OOmj2vXRoRbNq19F9VX4ix0sRt
w121Nd7sxybnx6n5YqiyG8m3k5vgihkb27yqjI5tM3av5hh14XY6UEO0u4zPdW42
OIahjmpolIR6G7BWI8gfVoQ/4f46totPCLCxxM99/INmmL9K1TVHNgXa9tisZrkp
HX0NlOhIsxkdCwAdBG/pwCzPLS2F4wjlKzCg97wrZEYoUVjcqE5eY0ixngVIynR4
LPlC0VS0wRFednJ8EvhK1Z6Q1bbjANCg7jfXsDDztadOV2wwaRGtLCsSjp16JMNT
XNDVoW9lv8jN+0UEETKC+MAm1/AMO6TrG3gRTK81Wue2LogzIxJd75jiIaL1QG9M
glkZ6vzi5uZYz2lVsE/E2c4PXjDMNHOLBK3eo4A+AGo+al/mh/fvEpBH8AW9qXRN
81EsGe3ls1NWsYzaNev6+bSVHs7WrGtgg2AUa9aZIcamO9Y1LptykjcHjiv06Z0C
WZTkPWRTpjnWuOdi6iCYXu88nBqE732/7HokQt6v8ws7f+isCID19TtNMV+Snw75
rxSQAHMmaigu90Z7V0FlbB1D7WYp4GAkGLiUilP+Xpje/4/U5PrgcB0G8qoOT5lE
ciH2BdicSAjROb+ws+Cl/iOVMrOm8lWq7Haczt6vSUDlNkeMIWLLhJChWEOfO5il
AKNtpp3VEUno21Izkb+fm8rI/++Qiug0hQLBG9jsqPxfNHPBp4WTmGBzauGyPHG9
C19fg1vnV+nA+rsiMfaroRlZ56pUuZvrC1CdSwkTJFbr43aQsvUJpnqOexP0XoDZ
SfsQ/DWUYsieL7UZagC0t09JTNq1ScNen9cPRdcgzq5wVVij697BtPJqCvQodU8D
QsQTx4mDKDcL2ZaXrrvuUo3qzvYbp7HN+uJRuMbLWSds1OoIEbeeAqf6mMHK525x
k58i+OxRBfHojxGPF9EGFPrzWsuidR0lZs6o21B0rLIxf6gCdSJISRMtWExiNPKb
gpzRn1nHefZFu7rokkMEHT1BYRW2x2LDYACpuvdpL4NI4vbUEstESBZOXGXAXSeV
Wk7Bf6J8dV89AtL/FPS4XWnRweR/RR2SZwFCbLvgngGOt7Vsri0Y/IdJiKCIDBgp
qM5MrMXRdKjsAIqmIX89vvcxMkcsm7bKvz47mxK/NO733pHPdAlDzd9onF7iTNjK
Ab/jQHvxo4E/AQrMFs+I/ZIfchNoh4/mFB2N2r6P2KwcIyAW9G2pve6557HSIzXs
hTy7OQweUrWbLguDJUGKA6vNSX1ncbYsPdpK0AbuWrIh/8WAgQ4lEd+RFS91G5fB
Mmb0krq3N/TmVK9Urt75rVxKYrBMP+Le8kEIJPRRhGpBAJyGcs1IptDaejzEjRg9
5Gaq1asXXbF9R3az0pcuw7nLAbE14dGXta7SJSkAnd9vqrg3HCzYJRRCF53Zyr+0
BmoyXQTLsVsz9jrYu5CnFy1wbOPNVCAaWhgyUs3OIS0rvFmHnrGVryIkyFsZvUPG
zxk/oSIrwF/DAZiLpVOCxa1p5LSk+6ryxdqLUshMWhviUMujsk4TdVsghJKM1C40
l5oZgcIDhkVAr30nBC+7xa1CHi46HHeQbaDYyyvZGDf6OWLvZ9XRernUsFvBwcl0
MR/K1cgfTqajR4xNpYhcJid3LUnQdfimZjOIe5uCWxuUalTG2vroedzKc77pgW9B
pPanzmkWq2o2/hMEX+zDofKxu+PD/7Ngq7EqURILtytKXs960F6/Hqf0cq6wUypt
3MiEOnCXNs62WM4q/yNspPdCYHVCsTdxXTXM1kguOov+vH2K558MCpDpCP+b5mfx
I/Zqv8dHaEH2PN2sjMKnR/TeKIy7kkz/mz/FBavlq74BIWO8oCHJJLjJEjhjjP7L
gBBtXRkqbrOlubzJAuuyJJHSqfN3nxJ+/oP+FsbQ/huhMS/y3qOmzUxIu5PqUfmR
DSo9UhA1uXmCqA9ZWWV/sOA/5+osYBTI7bNTs7no6DF9PLUzZbHKXTZD1pGj8UuS
IWdWHcROYpB1LnjqHRuQIgZW5YHE5ehT7a7LlvLpRvAT0qys4r6wDDIS4nn35ccp
nwjXNhKr9pKF5+50l8YERevEPl1Fv8pokIEPWIbwJK5TKXWY9It8VG/Z2yitVEta
QK2egAwvtR4VZLUzDkq/8Zms8HADOr2ltYkfHMuH0vIW1WOIngS82vxH1VYKsqHr
5tKmvlIwe0P+eyTn7ZYY7pXlT3ntBSjn5XkM7nFp9KhqPGXCr7TKPN5b6x+ICq5k
5l2MgnUBVj8hKL3ZcBq4Fr3/8lfdsRtonTeFNCQUQNBS8WTyEH5jAYrD/Ft2TnxO
KxEbBAjmAvHogml2MdCXadBbULLMsXXY0BVPHM8MDEbUHZ3SXWiANOxOh6f4V4Mw
bQBFkELfHRq9RvEH18oq/jrMuwUMv/tF23Yuh7wwF4HQ67FinobN/Nx1cfT/o3YD
AWTCVCv8LZc2tvmbHQpfXL517aoEDr7VAnG2F2ZXjJmObGw83T/UlB0z3kBFl9pI
hvpDb0+5dRx4hHetlI6K42VSbpdBdxQx3r1V1T2QX6NszGsdTiy/fOIV1RexNKpu
zvjVgffO/zHkrn/FOrWa5ONH/78Pxe6054mRku9CvYnO8+ggExE7p35WNbQhGY05
ZEn0lcLSiAgOVFZAKEqgScMNA+m0QNjkgBmUh/P0yikVmRAIfqddYRLRZjTwMuLw
ZK3GObs8xSADqh65Drzg79JrvBs/fDGpl8ThW87uXIiCuPpLxzwhD4VQD2EtLI9g
sxSPjCj8u4wFw6AFPSWymQ1dxGzICHZCX5gvxM6P8MSum/DUVOge6zbvMBI+6gF2
nphJ3XZGz8MsJG9MWGlhiitPtva6bNaxxJ2OBpCSVautQM6O7ptRJkFKVbBIU3xD
au6QZd+njXPMiKD2/B3X2qlp43xo/+J4A/OGL/sN8iu+bk1qyOV8Qva4CmfipliU
0jW6dmMNqMOcqiEMsNWNsn0Rh4Yh+qmAgHShpjEuzWhGYli1Y6WDtQbRiDkP4TFp
znP8mZN2dlQ+ghC7jb6Xdi5aRKwIbKvSV0sr/xHiJY+Bzq4SN2S7Ftfsi7RK8q5K
Gs5ELhwQY8i1jwmYgp63/duRYfvKskyG2aDtexZ2AtEXNhzymkSow5EFcpPWVj2b
CsAat9Mtv+IoWZvmvuHAIFRxeOEYpcx+yBEthEu0ZXxobsivps15z9cGUty9rzPE
Jh8GR6lsWxc06jpgKKlxptgrT0ClkMHuL+GA9/rlDGIs627XfWVey2RH4+In8Be3
987/7H7LF8IBfWy+T0xr3giDYErbhItcQtHk/m2X2lTLXj4fXx3FwEojh/10BEv6
2Ri5OZ3GNZTJND/98oVdk8+o/+132Y5jBEUyq9b8t7iuHYilhETxJjRhLSKlJxvp
g7O0CEr+QBB6ZOrk+Df6uHIMEofbvS0tL0zJWcptgFJbX1BSJ1DWpFa0X/2V5BJ2
GxzXp8p1qnSR6ZST/eq/O4D1GNGAXqhG7C6CWvzWu5X7zCczC9458QUSanY4VJ0L
g4eekGEeM/kESOM09XL9Z4paP3FY5nljiWOTiZnNxZqrV4ZrIfWeXvGICRd9WsSH
LuDJ6Pt5SRyYLBCYG0YMpu9ImizQe9Y+lbyIsUxw5oB3YjKHPdPcCvQ8nis0Hcxz
Pb+eTAdTBfG/X0ysQOWzz4GKCS5GDYD0fD5eV2Zuqav5tZjXTs4CgXDrwDqhvxDy
TEeYdH4SrwHiQb83nT2WTV8YgWnbdsgIv5GrRvgV9K06vBti+72sxvsDYkqyhHow
jqnnyBYahHHtoKwFtqCYqTViKK5I9d4oLLK+KC9oarEl3dcyKFUIvkc0ah+SUZYL
/H4BjB8P7JCMpJvAMoA+WSU/hUPwIrv9Wf2eHIJVUWl14SEXiUwU3V/cRBzeCPSX
ArZJNl1rO9i/eGjK0glVNKqJqW2OCsTxNQUslXLiZNwGgn2TXi+kU1fS/nFZkwP+
Gv7tLb1LlQSqLYBtEtlqu7Bq7KKqirq58MteLvB7q159I0uo5eEjBAa3EAtXEdab
v5k1hycAV2nMh39+yFHlD5eYV2mpoOASpTRy3X9UOjAtbQ2iiDr0ACY7PFwDob+c
cy2SmmISy+3qk6YwkDFNVNoFqcR5PHJi6lHh/UYqfB5Wzxz8/O45LTmoJltDVGJz
SmJo05EnPV56+0/LEVofQj/x40XIT6NYv4ShZoFdG3lSTAUeq7OJSGg3YC69IYf0
0CKi3fvous4/SNL5qUylZjOlViVa2Njav2XooGQVgX0W4Fz9s+RDgd5pClULPnwK
/uSIClpsrtNUhrZdFtZM2IOAHDawDj0L3l7iE/DwgWMm1xkeOuYg5Fge7q4zmPGd
6VsFGZDbNTnOglHLNxEDfRCPncNJhhj9OCLeKP/PWuLBjO+5sciTBDykYK+GMxkI
uIh9GKEcsVe9j/6CgxGLH5k7yk5nKY63mZ5Q3Fg+uo75nQi7ZDC3gEvZqMH1Ble3
0V8abz5v74IiUF1MjPPdJ0Rp3OUbHx21mLOsHMvDKU5kMcWLWjQSI+TjFB17fTLE
AC6dwiA2zRIn7PpCEEngcKIHfAtk9lz/194dbb8zOx6Ni53CPIp7x/yqmext+Xja
sR7ZaYS59be59gJz25IwnvARxjhVp17nNQRQPKh78x572ypbeJ+n2QPHCg1MOhLC
0FkB6E0CRc2+AklRxHiSt1JJ7KIkgRCNCDorrf010JPhBR/F/h+Rkew/JEbwTpUI
rDDBSAfshXzNgyw2nolpfGhjkqXszOUd+lhNleNs2FeGvdJyHxKrIQwc2xkEAKH4
3nYqHfQaq2hOb2HOojFZdOb3WE7hvEKCW3GxFeE26YYD6/MR8qlJ9aBCTe69wsAb
xy7WXf6/qf84BtHZfvXXDwgcNWB7vnny3CtiqnUXE9UF6HFmA+Pa3gazsMxKJDav
+gV3CJnvdn1la30G8UhGOXj0RzzfSwbsr40qKlv/F61M6zvknCztxCNVqTcwz2kP
67EHQRWJ9F+BUPIqur0jrreaawCgWy8gqpAolDogtaoaLKY1kfOQkWualf2RvWh4
eZO3VaLCNdZiY28aliF9XjGtFMPRnfoffJ1wQxT6luGuUh2nsq7g71b8G2uUgNVk
wvA3fTB4OrAYRtsWTaPK7ygPM/6xc01qfsDD77Y7KDCiUwTDBe3toagWfKflR7qT
SoEV+bghxIpSWAUKgI6xzzOC/H92LqKBQrbufXl0uwuSYuPSRuBDOnRtmNWofIGr
DK0BHzdLBepAKft7yo+6VYTy0Mb4VV3toZKlT9Mfw0PJh78GdSYj4iIelGivjWxE
hrRN3aLBH0t+/5c4uaqdkOFZsQGJ3iUAHtkIwye/9g2H47g/BgVcYW6CPfxrOQ6Y
WqTWR6mKpwm6XMbHCcKqDNEYfKZG/VFYkGXu9m2ABYauzjvIO1unba6PHp2A1wPh
+iD75yKQtcVnh6V2EqsTHS2M8pSXRyJRWo3xCF2ZY/mjyK/NepuBbCx/if32KVV1
MkuLQoduYm9tbqfplPukwATUfoFDFe8MKulHuiQGtoVGhQxs7KjUehILDZBPtEvy
Rbm5AFDEtZL0+eDM6WgyEn2R1FmzR/tJOKJmtf81aADdrQQJRBx4/s/aDLEcZIfj
jYfglxnFeKMTY6IwkuxcEacatG/akKCOcouFAIU9zEGs6ud3me4dmj78JFerN6pt
G6SHu9HA2ldJhCDKrIxDTP0wUH2ZBNsP9PRNBPjGRhYKD7yJ8z7J6+r/tex9axNE
zmPmzmBb8XjSLwrs1Pkhz/i/yfzglOzC2EPceasWexLJZmlp2EecnWiJTh9PiEhP
Z0PzPkFU0HynOkea8cI3kQWHL53DZjZ4/mok1gJ4yH5xsMbVJjEe45fMBZu7B4fM
A85ZosC+nj30zv8NJPMB/oDZHpMY2TjFwSoTbVhWGymWUAqvG6GLQNnyDTr7Wy7a
gNnMfwMsc+Og7f1O8ZK/ZOmBoz+k5xTHgkBYpQ0QLyrGhK/ex0UrFIb1q8pxeYf6
JWGcPtXOjmp0mfvUTKjcPk8RRm3wAQEOuRY6+4n+vbwX87Pe8knZc0916bKCTroy
hTWmLbKIWtD4rbG2gFs31hvPCOuhj+K16rIQoSnASN3EvOw6MMHkX5L4ssHCkZhO
McQ0OkGKjAektXFI07Yxlm8HQzSbB8Y/wuGrLtmS/HVG30x3YoT7WqQdFoAfdpBo
cICcFmLTYK16TzJt4KazSg2QZLoU5jrNiZWUE8AKRojlXMe5oCKSEQ2NrjsOYYFH
PJclmNoa4bbYkr/8bCVfSkXnhZV8zQjifQidOA7MisOFfm27rZedN7pu8a5bytb2
PRnkyNAKOVp3RyrA3aEy2xtBLXNJrBFl5zdIKNzqf2wC4vx5dEUOKP+4cl6j2Kdq
vDgyxfdOXUIuueRbSfVZr7Ld9h45bVXU8oYdbWpfLqqkNjeEz/cxTOWju+ktg73P
NiOhw8DgCkz7u6hAqkK6c0E95kgn1n7RIJLa7ubIInATequlYQkaULc8VtDBR4iE
UQwJGF926VQKkJ0QeJuLE6Vbmgivfw920B0M3wQJx4IeX8LslVNYj6Iq1lpxls/T
WzsxGM4KMbtn9YCrykfsMLnZYowuDv19GJyDNZuR2Oj404O7OdB+SZMshBEzVak3
j6nQ0Gc+ymxjlkO2jKI3BigX7jNx4lnK7p5j+kvbS1xZRgTaC2QgBdy+ZEzleh7i
rvuws6de9xuLVT9oOaSf7jNO/7CDtiJfKc/wimUEozCb95/hJqrDuEHHiQNZr7cM
OKSd5GdR/Ky2elqyN7xXckM7EgwDv9GXG5mGUvf6egBIaZJwOyGO6V4kyweOaHSy
I9HQNv0nfSZw1YmQqP71i2nkJostW/bf30h+lqfp7Yln/aF4QBv0TzH2kX+bQQ6S
oHuCQRzWQlnBz9BvtbsShU7PX6kX8erd/bU1jI0o5ZZuF95S+17UxoRqnZ3Odgta
9L1sAa8ciz0gnyZYL4wyhDBrPKQgxEP3b+7s2ybFQNfVgJS8UY+hY7ksZTqE5D1D
UOIgZ5o2e4XTk5IzWOXos78kWkDcM2l64z41lfU3mUUykv4wup8r3ROWNwadDuva
RNqTkrhzLyU4ovf0gD+E5FHPTBygTv7H1wWqAIWMKQgl1QdU7w6LSLFKszucrJIl
vHFQnB83Q1t0g0/TPKuqU/cyIvSzw52ePYlbz1f3ppoQUgozI/1zoXoT05yKJQ5b
SNCly8ZlLT/FDN4sBAYDzfifqbKl5MoAoLG6+eShTroEDjT8CEmcTystk6t3Duu6
tWzjhU8s0auL/MKC9lyu0h5qav5/HgSTeZZhK6LpaZ8Uxnqneyll82HVKtsPUkgD
E/AUTW/qGyJatUVB8xynvcSxlfMC/EXtzzK+NlqVWZcHj9cbBH8BkDiRSbHfN1xC
RtzoZimhTZBTJOvJg0w7l0D0rEValJ2xQYi8vuQ/0bWkjpmMmvK0AyMa+wepXb2F
9ZIEg6B/5wr8r8g42xtfa1PLdiTZqHURrTRncV8oTI4DvZMSctaXgXlhNS5FpUor
Gy7Pr9cbLVT7738TBDCSHaAvymj4MWkq1oifhpkO8XmLouOrbWV/F6vJzPTnZn7m
OPpWAmSPCAt9I+OUBiEkKs0o5MuwzJ0U/yZEtlFsTz633vf+eY00FqpeCrQ0+ClR
jqKdudRKTuqxbp+pJc5MKc1AsrfX+qiwExzTFqr6DovBFQHFwxRyeZjwh6wjk0a3

//pragma protect end_data_block
//pragma protect digest_block
BbsHfjV9RZjwwm0xeDyWwttIJ8g=
//pragma protect end_digest_block
//pragma protect end_protected
